module Motion_Update_input_selector
#(
	parameter DATA_WIDTH									= 32,
	parameter GLOBAL_CELL_ADDR_LEN					= 7,
	parameter TOTAL_CELL_NUM							= 64
)
(
	input clk,
	input rst,
	input [GLOBAL_CELL_ADDR_LEN-1:0] cell_being_updated_id, 
	input [TOTAL_CELL_NUM*3*DATA_WIDTH-1:0] all_Motion_Update_velocity_data,
	input [TOTAL_CELL_NUM*3*DATA_WIDTH-1:0] all_Motion_Update_position_data,
	input [TOTAL_CELL_NUM*3*DATA_WIDTH-1:0] all_Motion_Update_force_data,
	input Motion_Update_enable,
	
	output [TOTAL_CELL_NUM-1:0] motion_update_to_cache_read_force_request,
	output [3*DATA_WIDTH-1:0] Motion_Update_velocity_data,
	output [3*DATA_WIDTH-1:0] Motion_Update_position_data,
	output [3*DATA_WIDTH-1:0] Motion_Update_force_data
);

reg [3*DATA_WIDTH-1:0] reg_Motion_Update_velocity_data;
reg [3*DATA_WIDTH-1:0] reg_Motion_Update_position_data;
reg [3*DATA_WIDTH-1:0] reg_Motion_Update_force_data;
reg [TOTAL_CELL_NUM-1:0] reg_motion_update_to_cache_read_force_request;
assign Motion_Update_velocity_data = reg_Motion_Update_velocity_data;
assign Motion_Update_position_data = reg_Motion_Update_position_data;
assign Motion_Update_force_data = reg_Motion_Update_force_data;
assign motion_update_to_cache_read_force_request = reg_motion_update_to_cache_read_force_request;
	
always@(*)
	begin
	if (rst)
		begin
		reg_motion_update_to_cache_read_force_request <= 0;
		reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= 0;
		reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= 0;
		reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= 0;
		end
	else
		begin
		reg_motion_update_to_cache_read_force_request <= Motion_Update_enable << (cell_being_updated_id-1);
		case(cell_being_updated_id)
			1:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH];
				end
			2:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH];
				end
			3:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH];
				end
			4:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH];
				end
			5:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH];
				end
			6:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH];
				end
			7:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH];
				end
			8:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH];
				end
			9:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[9*3*DATA_WIDTH-1:8*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[9*3*DATA_WIDTH-1:8*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[9*3*DATA_WIDTH-1:8*3*DATA_WIDTH];
				end
			10:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[10*3*DATA_WIDTH-1:9*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[10*3*DATA_WIDTH-1:9*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[10*3*DATA_WIDTH-1:9*3*DATA_WIDTH];
				end
			11:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[11*3*DATA_WIDTH-1:10*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[11*3*DATA_WIDTH-1:10*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[11*3*DATA_WIDTH-1:10*3*DATA_WIDTH];
				end
			12:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[12*3*DATA_WIDTH-1:11*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[12*3*DATA_WIDTH-1:11*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[12*3*DATA_WIDTH-1:11*3*DATA_WIDTH];
				end
			13:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[13*3*DATA_WIDTH-1:12*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[13*3*DATA_WIDTH-1:12*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[13*3*DATA_WIDTH-1:12*3*DATA_WIDTH];
				end
			14:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[14*3*DATA_WIDTH-1:13*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[14*3*DATA_WIDTH-1:13*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[14*3*DATA_WIDTH-1:13*3*DATA_WIDTH];
				end
			15:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[15*3*DATA_WIDTH-1:14*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[15*3*DATA_WIDTH-1:14*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[15*3*DATA_WIDTH-1:14*3*DATA_WIDTH];
				end
			16:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[16*3*DATA_WIDTH-1:15*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[16*3*DATA_WIDTH-1:15*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[16*3*DATA_WIDTH-1:15*3*DATA_WIDTH];
				end
			17:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH];
				end
			18:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH];
				end
			19:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH];
				end
			20:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH];
				end
			21:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH];
				end
			22:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH];
				end
			23:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH];
				end
			24:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH];
				end
			25:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[25*3*DATA_WIDTH-1:24*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[25*3*DATA_WIDTH-1:24*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[25*3*DATA_WIDTH-1:24*3*DATA_WIDTH];
				end
			26:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[26*3*DATA_WIDTH-1:25*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[26*3*DATA_WIDTH-1:25*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[26*3*DATA_WIDTH-1:25*3*DATA_WIDTH];
				end
			27:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[27*3*DATA_WIDTH-1:26*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[27*3*DATA_WIDTH-1:26*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[27*3*DATA_WIDTH-1:26*3*DATA_WIDTH];
				end
			28:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[28*3*DATA_WIDTH-1:27*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[28*3*DATA_WIDTH-1:27*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[28*3*DATA_WIDTH-1:27*3*DATA_WIDTH];
				end
			29:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH];
				end
			30:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH];
				end
			31:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH];
				end
			32:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH];
				end
			33:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[33*3*DATA_WIDTH-1:32*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[33*3*DATA_WIDTH-1:32*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[33*3*DATA_WIDTH-1:32*3*DATA_WIDTH];
				end
			34:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[34*3*DATA_WIDTH-1:33*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[34*3*DATA_WIDTH-1:33*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[34*3*DATA_WIDTH-1:33*3*DATA_WIDTH];
				end
			35:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[35*3*DATA_WIDTH-1:34*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[35*3*DATA_WIDTH-1:34*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[35*3*DATA_WIDTH-1:34*3*DATA_WIDTH];
				end
			36:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[36*3*DATA_WIDTH-1:35*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[36*3*DATA_WIDTH-1:35*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[36*3*DATA_WIDTH-1:35*3*DATA_WIDTH];
				end
			37:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[37*3*DATA_WIDTH-1:36*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[37*3*DATA_WIDTH-1:36*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[37*3*DATA_WIDTH-1:36*3*DATA_WIDTH];
				end
			38:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[38*3*DATA_WIDTH-1:37*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[38*3*DATA_WIDTH-1:37*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[38*3*DATA_WIDTH-1:37*3*DATA_WIDTH];
				end
			39:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[39*3*DATA_WIDTH-1:38*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[39*3*DATA_WIDTH-1:38*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[39*3*DATA_WIDTH-1:38*3*DATA_WIDTH];
				end
			40:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[40*3*DATA_WIDTH-1:39*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[40*3*DATA_WIDTH-1:39*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[40*3*DATA_WIDTH-1:39*3*DATA_WIDTH];
				end
			41:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[41*3*DATA_WIDTH-1:40*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[41*3*DATA_WIDTH-1:40*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[41*3*DATA_WIDTH-1:40*3*DATA_WIDTH];
				end
			42:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[42*3*DATA_WIDTH-1:41*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[42*3*DATA_WIDTH-1:41*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[42*3*DATA_WIDTH-1:41*3*DATA_WIDTH];
				end
			43:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[43*3*DATA_WIDTH-1:42*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[43*3*DATA_WIDTH-1:42*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[43*3*DATA_WIDTH-1:42*3*DATA_WIDTH];
				end
			44:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[44*3*DATA_WIDTH-1:43*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[44*3*DATA_WIDTH-1:43*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[44*3*DATA_WIDTH-1:43*3*DATA_WIDTH];
				end
			45:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[45*3*DATA_WIDTH-1:44*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[45*3*DATA_WIDTH-1:44*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[45*3*DATA_WIDTH-1:44*3*DATA_WIDTH];
				end
			46:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[46*3*DATA_WIDTH-1:45*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[46*3*DATA_WIDTH-1:45*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[46*3*DATA_WIDTH-1:45*3*DATA_WIDTH];
				end
			47:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[47*3*DATA_WIDTH-1:46*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[47*3*DATA_WIDTH-1:46*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[47*3*DATA_WIDTH-1:46*3*DATA_WIDTH];
				end
			48:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[48*3*DATA_WIDTH-1:47*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[48*3*DATA_WIDTH-1:47*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[48*3*DATA_WIDTH-1:47*3*DATA_WIDTH];
				end
			49:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[49*3*DATA_WIDTH-1:48*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[49*3*DATA_WIDTH-1:48*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[49*3*DATA_WIDTH-1:48*3*DATA_WIDTH];
				end
			50:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[50*3*DATA_WIDTH-1:49*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[50*3*DATA_WIDTH-1:49*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[50*3*DATA_WIDTH-1:49*3*DATA_WIDTH];
				end
			51:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[51*3*DATA_WIDTH-1:50*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[51*3*DATA_WIDTH-1:50*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[51*3*DATA_WIDTH-1:50*3*DATA_WIDTH];
				end
			52:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[52*3*DATA_WIDTH-1:51*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[52*3*DATA_WIDTH-1:51*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[52*3*DATA_WIDTH-1:51*3*DATA_WIDTH];
				end
			53:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[53*3*DATA_WIDTH-1:52*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[53*3*DATA_WIDTH-1:52*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[53*3*DATA_WIDTH-1:52*3*DATA_WIDTH];
				end
			54:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[54*3*DATA_WIDTH-1:53*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[54*3*DATA_WIDTH-1:53*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[54*3*DATA_WIDTH-1:53*3*DATA_WIDTH];
				end
			55:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[55*3*DATA_WIDTH-1:54*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[55*3*DATA_WIDTH-1:54*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[55*3*DATA_WIDTH-1:54*3*DATA_WIDTH];
				end
			56:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[56*3*DATA_WIDTH-1:55*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[56*3*DATA_WIDTH-1:55*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[56*3*DATA_WIDTH-1:55*3*DATA_WIDTH];
				end
			57:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[57*3*DATA_WIDTH-1:56*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[57*3*DATA_WIDTH-1:56*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[57*3*DATA_WIDTH-1:56*3*DATA_WIDTH];
				end
			58:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[58*3*DATA_WIDTH-1:57*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[58*3*DATA_WIDTH-1:57*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[58*3*DATA_WIDTH-1:57*3*DATA_WIDTH];
				end
			59:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[59*3*DATA_WIDTH-1:58*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[59*3*DATA_WIDTH-1:58*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[59*3*DATA_WIDTH-1:58*3*DATA_WIDTH];
				end
			60:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[60*3*DATA_WIDTH-1:59*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[60*3*DATA_WIDTH-1:59*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[60*3*DATA_WIDTH-1:59*3*DATA_WIDTH];
				end
			61:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[61*3*DATA_WIDTH-1:60*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[61*3*DATA_WIDTH-1:60*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[61*3*DATA_WIDTH-1:60*3*DATA_WIDTH];
				end
			62:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[62*3*DATA_WIDTH-1:61*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[62*3*DATA_WIDTH-1:61*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[62*3*DATA_WIDTH-1:61*3*DATA_WIDTH];
				end
			63:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[63*3*DATA_WIDTH-1:62*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[63*3*DATA_WIDTH-1:62*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[63*3*DATA_WIDTH-1:62*3*DATA_WIDTH];
				end
			64:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_velocity_data[64*3*DATA_WIDTH-1:63*3*DATA_WIDTH];
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_position_data[64*3*DATA_WIDTH-1:63*3*DATA_WIDTH];
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= all_Motion_Update_force_data[64*3*DATA_WIDTH-1:63*3*DATA_WIDTH];
				end
			default:
				begin
				reg_Motion_Update_velocity_data[3*DATA_WIDTH-1:0] <= 0;
				reg_Motion_Update_position_data[3*DATA_WIDTH-1:0] <= 0;
				reg_Motion_Update_force_data[3*DATA_WIDTH-1:0] <= 0;
				end
		endcase
		end
	end

endmodule