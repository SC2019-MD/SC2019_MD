/*****************************************************
Used to store all the position caches, nice and clean
*****************************************************/
module All_Position_Caches_64_Cells
#(
	parameter DATA_WIDTH 					= 32,
	parameter CELL_ID_WIDTH					= 4,
	parameter TOTAL_CELL_NUM				= 64,
	parameter MAX_CELL_PARTICLE_NUM		= 100,
	parameter CELL_ADDR_WIDTH				= 7
)
(
	input clk,
	input rst,
	input Motion_Update_enable,
	input [CELL_ADDR_WIDTH-1:0] Motion_Update_position_read_addr,
	input [TOTAL_CELL_NUM*CELL_ADDR_WIDTH-1:0] FSM_to_Cell_read_addr,
	input [3*DATA_WIDTH-1:0] Motion_Update_out_position_data,
	input [3*CELL_ID_WIDTH-1:0] Motion_Update_dst_cell,
	input Motion_Update_out_position_data_valid,
	input Motion_Update_position_read_en,
	input [TOTAL_CELL_NUM-1:0] FSM_to_Cell_rden,
	
	output [TOTAL_CELL_NUM*3*DATA_WIDTH-1:0] Position_Cache_readout_position
);
		
	Pos_Cache_1_1_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(1)
	)
	cell_1_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[0]),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_1_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(2)
	)
	cell_1_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[1]),
		.out_particle_info(Position_Cache_readout_position[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_1_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(3)
	)
	cell_1_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[2]),
		.out_particle_info(Position_Cache_readout_position[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_1_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(4)
	)
	cell_1_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[3]),
		.out_particle_info(Position_Cache_readout_position[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_2_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(1)
	)
	cell_1_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[4]),
		.out_particle_info(Position_Cache_readout_position[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(2)
	)
	cell_1_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[5]),
		.out_particle_info(Position_Cache_readout_position[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_2_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(3)
	)
	cell_1_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[6]),
		.out_particle_info(Position_Cache_readout_position[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_2_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(4)
	)
	cell_1_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[7]),
		.out_particle_info(Position_Cache_readout_position[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_3_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(1)
	)
	cell_1_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[8]),
		.out_particle_info(Position_Cache_readout_position[9*3*DATA_WIDTH-1:8*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_3_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(2)
	)
	cell_1_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[9]),
		.out_particle_info(Position_Cache_readout_position[10*3*DATA_WIDTH-1:9*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_3_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(3)
	)
	cell_1_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[10]),
		.out_particle_info(Position_Cache_readout_position[11*3*DATA_WIDTH-1:10*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_3_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(4)
	)
	cell_1_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[11]),
		.out_particle_info(Position_Cache_readout_position[12*3*DATA_WIDTH-1:11*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_4_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(1)
	)
	cell_1_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[12]),
		.out_particle_info(Position_Cache_readout_position[13*3*DATA_WIDTH-1:12*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_4_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(2)
	)
	cell_1_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[13]),
		.out_particle_info(Position_Cache_readout_position[14*3*DATA_WIDTH-1:13*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_4_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(3)
	)
	cell_1_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[15*CELL_ADDR_WIDTH-1:14*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[14]),
		.out_particle_info(Position_Cache_readout_position[15*3*DATA_WIDTH-1:14*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_4_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(4)
	)
	cell_1_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[16*CELL_ADDR_WIDTH-1:15*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[15]),
		.out_particle_info(Position_Cache_readout_position[16*3*DATA_WIDTH-1:15*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_1_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(1)
	)
	cell_2_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[17*CELL_ADDR_WIDTH-1:16*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[16]),
		.out_particle_info(Position_Cache_readout_position[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_1_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(2)
	)
	cell_2_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[18*CELL_ADDR_WIDTH-1:17*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[17]),
		.out_particle_info(Position_Cache_readout_position[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_1_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(3)
	)
	cell_2_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[19*CELL_ADDR_WIDTH-1:18*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[18]),
		.out_particle_info(Position_Cache_readout_position[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_1_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(4)
	)
	cell_2_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[20*CELL_ADDR_WIDTH-1:19*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[19]),
		.out_particle_info(Position_Cache_readout_position[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_2_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(1)
	)
	cell_2_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[21*CELL_ADDR_WIDTH-1:20*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[20]),
		.out_particle_info(Position_Cache_readout_position[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(2)
	)
	cell_2_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[22*CELL_ADDR_WIDTH-1:21*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[21]),
		.out_particle_info(Position_Cache_readout_position[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_2_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(3)
	)
	cell_2_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[23*CELL_ADDR_WIDTH-1:22*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[22]),
		.out_particle_info(Position_Cache_readout_position[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_2_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(4)
	)
	cell_2_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[24*CELL_ADDR_WIDTH-1:23*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[23]),
		.out_particle_info(Position_Cache_readout_position[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_3_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(1)
	)
	cell_2_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[25*CELL_ADDR_WIDTH-1:24*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[24]),
		.out_particle_info(Position_Cache_readout_position[25*3*DATA_WIDTH-1:24*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_3_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(2)
	)
	cell_2_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[26*CELL_ADDR_WIDTH-1:25*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[25]),
		.out_particle_info(Position_Cache_readout_position[26*3*DATA_WIDTH-1:25*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_3_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(3)
	)
	cell_2_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[27*CELL_ADDR_WIDTH-1:26*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[26]),
		.out_particle_info(Position_Cache_readout_position[27*3*DATA_WIDTH-1:26*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_3_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(4)
	)
	cell_2_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[28*CELL_ADDR_WIDTH-1:27*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[27]),
		.out_particle_info(Position_Cache_readout_position[28*3*DATA_WIDTH-1:27*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_4_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(1)
	)
	cell_2_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[29*CELL_ADDR_WIDTH-1:28*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[28]),
		.out_particle_info(Position_Cache_readout_position[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_4_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(2)
	)
	cell_2_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[30*CELL_ADDR_WIDTH-1:29*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[29]),
		.out_particle_info(Position_Cache_readout_position[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_4_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(3)
	)
	cell_2_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[31*CELL_ADDR_WIDTH-1:30*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[30]),
		.out_particle_info(Position_Cache_readout_position[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_4_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(4)
	)
	cell_2_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[32*CELL_ADDR_WIDTH-1:31*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[31]),
		.out_particle_info(Position_Cache_readout_position[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_1_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(1)
	)
	cell_3_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[33*CELL_ADDR_WIDTH-1:32*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[32]),
		.out_particle_info(Position_Cache_readout_position[33*3*DATA_WIDTH-1:32*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_1_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(2)
	)
	cell_3_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[34*CELL_ADDR_WIDTH-1:33*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[33]),
		.out_particle_info(Position_Cache_readout_position[34*3*DATA_WIDTH-1:33*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_1_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(3)
	)
	cell_3_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[35*CELL_ADDR_WIDTH-1:34*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[34]),
		.out_particle_info(Position_Cache_readout_position[35*3*DATA_WIDTH-1:34*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_1_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(4)
	)
	cell_3_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[36*CELL_ADDR_WIDTH-1:35*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[35]),
		.out_particle_info(Position_Cache_readout_position[36*3*DATA_WIDTH-1:35*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_2_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(1)
	)
	cell_3_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[37*CELL_ADDR_WIDTH-1:36*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[36]),
		.out_particle_info(Position_Cache_readout_position[37*3*DATA_WIDTH-1:36*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(2)
	)
	cell_3_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[38*CELL_ADDR_WIDTH-1:37*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[37]),
		.out_particle_info(Position_Cache_readout_position[38*3*DATA_WIDTH-1:37*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_2_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(3)
	)
	cell_3_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[39*CELL_ADDR_WIDTH-1:38*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[38]),
		.out_particle_info(Position_Cache_readout_position[39*3*DATA_WIDTH-1:38*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_2_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(4)
	)
	cell_3_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[40*CELL_ADDR_WIDTH-1:39*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[39]),
		.out_particle_info(Position_Cache_readout_position[40*3*DATA_WIDTH-1:39*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_3_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(1)
	)
	cell_3_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[41*CELL_ADDR_WIDTH-1:40*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[40]),
		.out_particle_info(Position_Cache_readout_position[41*3*DATA_WIDTH-1:40*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_3_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(2)
	)
	cell_3_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[42*CELL_ADDR_WIDTH-1:41*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[41]),
		.out_particle_info(Position_Cache_readout_position[42*3*DATA_WIDTH-1:41*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_3_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(3)
	)
	cell_3_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[43*CELL_ADDR_WIDTH-1:42*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[42]),
		.out_particle_info(Position_Cache_readout_position[43*3*DATA_WIDTH-1:42*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_3_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(4)
	)
	cell_3_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[44*CELL_ADDR_WIDTH-1:43*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[43]),
		.out_particle_info(Position_Cache_readout_position[44*3*DATA_WIDTH-1:43*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_4_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(1)
	)
	cell_3_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[45*CELL_ADDR_WIDTH-1:44*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[44]),
		.out_particle_info(Position_Cache_readout_position[45*3*DATA_WIDTH-1:44*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_4_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(2)
	)
	cell_3_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[46*CELL_ADDR_WIDTH-1:45*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[45]),
		.out_particle_info(Position_Cache_readout_position[46*3*DATA_WIDTH-1:45*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_4_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(3)
	)
	cell_3_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[47*CELL_ADDR_WIDTH-1:46*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[46]),
		.out_particle_info(Position_Cache_readout_position[47*3*DATA_WIDTH-1:46*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_4_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(4)
	)
	cell_3_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[48*CELL_ADDR_WIDTH-1:47*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[47]),
		.out_particle_info(Position_Cache_readout_position[48*3*DATA_WIDTH-1:47*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_1_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(1)
	)
	cell_4_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[49*CELL_ADDR_WIDTH-1:48*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[48]),
		.out_particle_info(Position_Cache_readout_position[49*3*DATA_WIDTH-1:48*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_1_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(2)
	)
	cell_4_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[50*CELL_ADDR_WIDTH-1:49*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[49]),
		.out_particle_info(Position_Cache_readout_position[50*3*DATA_WIDTH-1:49*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_1_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(3)
	)
	cell_4_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[51*CELL_ADDR_WIDTH-1:50*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[50]),
		.out_particle_info(Position_Cache_readout_position[51*3*DATA_WIDTH-1:50*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_1_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(4)
	)
	cell_4_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[52*CELL_ADDR_WIDTH-1:51*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[51]),
		.out_particle_info(Position_Cache_readout_position[52*3*DATA_WIDTH-1:51*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_2_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(1)
	)
	cell_4_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[53*CELL_ADDR_WIDTH-1:52*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[52]),
		.out_particle_info(Position_Cache_readout_position[53*3*DATA_WIDTH-1:52*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(2)
	)
	cell_4_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[54*CELL_ADDR_WIDTH-1:53*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[53]),
		.out_particle_info(Position_Cache_readout_position[54*3*DATA_WIDTH-1:53*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_2_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(3)
	)
	cell_4_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[55*CELL_ADDR_WIDTH-1:54*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[54]),
		.out_particle_info(Position_Cache_readout_position[55*3*DATA_WIDTH-1:54*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_2_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(4)
	)
	cell_4_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[56*CELL_ADDR_WIDTH-1:55*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[55]),
		.out_particle_info(Position_Cache_readout_position[56*3*DATA_WIDTH-1:55*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_3_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(1)
	)
	cell_4_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[57*CELL_ADDR_WIDTH-1:56*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[56]),
		.out_particle_info(Position_Cache_readout_position[57*3*DATA_WIDTH-1:56*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_3_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(2)
	)
	cell_4_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[58*CELL_ADDR_WIDTH-1:57*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[57]),
		.out_particle_info(Position_Cache_readout_position[58*3*DATA_WIDTH-1:57*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_3_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(3)
	)
	cell_4_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[59*CELL_ADDR_WIDTH-1:58*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[58]),
		.out_particle_info(Position_Cache_readout_position[59*3*DATA_WIDTH-1:58*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_3_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(4)
	)
	cell_4_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[60*CELL_ADDR_WIDTH-1:59*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[59]),
		.out_particle_info(Position_Cache_readout_position[60*3*DATA_WIDTH-1:59*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_4_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(1)
	)
	cell_4_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[61*CELL_ADDR_WIDTH-1:60*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[60]),
		.out_particle_info(Position_Cache_readout_position[61*3*DATA_WIDTH-1:60*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_4_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(2)
	)
	cell_4_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[62*CELL_ADDR_WIDTH-1:61*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[61]),
		.out_particle_info(Position_Cache_readout_position[62*3*DATA_WIDTH-1:61*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_4_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(3)
	)
	cell_4_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[63*CELL_ADDR_WIDTH-1:62*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[62]),
		.out_particle_info(Position_Cache_readout_position[63*3*DATA_WIDTH-1:62*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_4_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(4)
	)
	cell_4_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[64*CELL_ADDR_WIDTH-1:63*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden[63]),
		.out_particle_info(Position_Cache_readout_position[64*3*DATA_WIDTH-1:63*3*DATA_WIDTH])
	);
	
endmodule