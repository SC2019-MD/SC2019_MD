/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Module: fp_div.v
//
//	Function:
//				Wrapper on top of FP_DIV, to meet the port configuration in the old design
//
// Dependency:
//				FP_DIV.v
//
// Latency: 38 cycles
//
//
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module fp_div
#(
	parameter DATA_WIDTH = 32
)
(
	input clk,
	input [DATA_WIDTH-1:0] in1,
	input [DATA_WIDTH-1:0] in2,
	output [DATA_WIDTH-1:0] result
);

	FP_DIV FP_DIV
	(
		.clk(clk),
		.areset(1'b0),
		.a(in1),
		.b(in2),
		.q(result)
	);

endmodule
