/*****************************************************
Used to store all the velocity caches, nice and clean
*****************************************************/
module All_Velocity_Caches_64_Cells
#(
	parameter DATA_WIDTH 					= 32,
	parameter CELL_ID_WIDTH					= 4,
	parameter TOTAL_CELL_NUM				= 64,
	parameter MAX_CELL_PARTICLE_NUM		= 290,
	parameter CELL_ADDR_WIDTH				= 9
)
(
	input clk,
	input rst,
	input Motion_Update_enable,
	input [CELL_ADDR_WIDTH-1:0] Motion_Update_velocity_read_addr,
	input [3*DATA_WIDTH-1:0] Motion_Update_out_velocity_data,
	input [3*CELL_ID_WIDTH-1:0] Motion_Update_dst_cell,
	input Motion_Update_out_velocity_data_valid,
	input Motion_Update_velocity_read_en,
	
	output [TOTAL_CELL_NUM*3*DATA_WIDTH-1:0] Motion_Update_velocity_data
);


	Velocity_Cache_1_1_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd1),
		.CELL_Y(4'd1),
		.CELL_Z(4'd1)
	)
	Velocity_Cache_1_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	);
	Velocity_Cache_1_1_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd1),
		.CELL_Y(4'd1),
		.CELL_Z(4'd2)
	)
	Velocity_Cache_1_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH])
	);
	Velocity_Cache_1_1_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd1),
		.CELL_Y(4'd1),
		.CELL_Z(4'd3)
	)
	Velocity_Cache_1_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH])
	);
	Velocity_Cache_1_1_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd1),
		.CELL_Y(4'd1),
		.CELL_Z(4'd4)
	)
	Velocity_Cache_1_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH])
	);
	Velocity_Cache_1_2_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd1),
		.CELL_Y(4'd2),
		.CELL_Z(4'd1)
	)
	Velocity_Cache_1_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH])
	);
	Velocity_Cache_1_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd1),
		.CELL_Y(4'd2),
		.CELL_Z(4'd2)
	)
	Velocity_Cache_1_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH])
	);
	Velocity_Cache_1_2_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd1),
		.CELL_Y(4'd2),
		.CELL_Z(4'd3)
	)
	Velocity_Cache_1_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH])
	);
	Velocity_Cache_1_2_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd1),
		.CELL_Y(4'd2),
		.CELL_Z(4'd4)
	)
	Velocity_Cache_1_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH])
	);
	Velocity_Cache_1_3_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd1),
		.CELL_Y(4'd3),
		.CELL_Z(4'd1)
	)
	Velocity_Cache_1_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[9*3*DATA_WIDTH-1:8*3*DATA_WIDTH])
	);
	Velocity_Cache_1_3_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd1),
		.CELL_Y(4'd3),
		.CELL_Z(4'd2)
	)
	Velocity_Cache_1_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[10*3*DATA_WIDTH-1:9*3*DATA_WIDTH])
	);
	Velocity_Cache_1_3_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd1),
		.CELL_Y(4'd3),
		.CELL_Z(4'd3)
	)
	Velocity_Cache_1_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[11*3*DATA_WIDTH-1:10*3*DATA_WIDTH])
	);
	Velocity_Cache_1_3_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd1),
		.CELL_Y(4'd3),
		.CELL_Z(4'd4)
	)
	Velocity_Cache_1_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[12*3*DATA_WIDTH-1:11*3*DATA_WIDTH])
	);
	Velocity_Cache_1_4_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd1),
		.CELL_Y(4'd4),
		.CELL_Z(4'd1)
	)
	Velocity_Cache_1_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[13*3*DATA_WIDTH-1:12*3*DATA_WIDTH])
	);
	Velocity_Cache_1_4_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd1),
		.CELL_Y(4'd4),
		.CELL_Z(4'd2)
	)
	Velocity_Cache_1_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[14*3*DATA_WIDTH-1:13*3*DATA_WIDTH])
	);
	Velocity_Cache_1_4_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd1),
		.CELL_Y(4'd4),
		.CELL_Z(4'd3)
	)
	Velocity_Cache_1_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[15*3*DATA_WIDTH-1:14*3*DATA_WIDTH])
	);
	Velocity_Cache_1_4_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd1),
		.CELL_Y(4'd4),
		.CELL_Z(4'd4)
	)
	Velocity_Cache_1_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[16*3*DATA_WIDTH-1:15*3*DATA_WIDTH])
	);
	Velocity_Cache_2_1_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd2),
		.CELL_Y(4'd1),
		.CELL_Z(4'd1)
	)
	Velocity_Cache_2_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH])
	);
	Velocity_Cache_2_1_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd2),
		.CELL_Y(4'd1),
		.CELL_Z(4'd2)
	)
	Velocity_Cache_2_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH])
	);
	Velocity_Cache_2_1_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd2),
		.CELL_Y(4'd1),
		.CELL_Z(4'd3)
	)
	Velocity_Cache_2_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH])
	);
	Velocity_Cache_2_1_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd2),
		.CELL_Y(4'd1),
		.CELL_Z(4'd4)
	)
	Velocity_Cache_2_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH])
	);
	Velocity_Cache_2_2_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd2),
		.CELL_Y(4'd2),
		.CELL_Z(4'd1)
	)
	Velocity_Cache_2_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH])
	);
	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd2),
		.CELL_Y(4'd2),
		.CELL_Z(4'd2)
	)
	Velocity_Cache_2_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH])
	);
	Velocity_Cache_2_2_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd2),
		.CELL_Y(4'd2),
		.CELL_Z(4'd3)
	)
	Velocity_Cache_2_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH])
	);
	Velocity_Cache_2_2_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd2),
		.CELL_Y(4'd2),
		.CELL_Z(4'd4)
	)
	Velocity_Cache_2_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH])
	);
	Velocity_Cache_2_3_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd2),
		.CELL_Y(4'd3),
		.CELL_Z(4'd1)
	)
	Velocity_Cache_2_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[25*3*DATA_WIDTH-1:24*3*DATA_WIDTH])
	);
	Velocity_Cache_2_3_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd2),
		.CELL_Y(4'd3),
		.CELL_Z(4'd2)
	)
	Velocity_Cache_2_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[26*3*DATA_WIDTH-1:25*3*DATA_WIDTH])
	);
	Velocity_Cache_2_3_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd2),
		.CELL_Y(4'd3),
		.CELL_Z(4'd3)
	)
	Velocity_Cache_2_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[27*3*DATA_WIDTH-1:26*3*DATA_WIDTH])
	);
	Velocity_Cache_2_3_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd2),
		.CELL_Y(4'd3),
		.CELL_Z(4'd4)
	)
	Velocity_Cache_2_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[28*3*DATA_WIDTH-1:27*3*DATA_WIDTH])
	);
	Velocity_Cache_2_4_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd2),
		.CELL_Y(4'd4),
		.CELL_Z(4'd1)
	)
	Velocity_Cache_2_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH])
	);
	Velocity_Cache_2_4_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd2),
		.CELL_Y(4'd4),
		.CELL_Z(4'd2)
	)
	Velocity_Cache_2_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH])
	);
	Velocity_Cache_2_4_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd2),
		.CELL_Y(4'd4),
		.CELL_Z(4'd3)
	)
	Velocity_Cache_2_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH])
	);
	Velocity_Cache_2_4_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd2),
		.CELL_Y(4'd4),
		.CELL_Z(4'd4)
	)
	Velocity_Cache_2_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH])
	);
	Velocity_Cache_3_1_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd3),
		.CELL_Y(4'd1),
		.CELL_Z(4'd1)
	)
	Velocity_Cache_3_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[33*3*DATA_WIDTH-1:32*3*DATA_WIDTH])
	);
	Velocity_Cache_3_1_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd3),
		.CELL_Y(4'd1),
		.CELL_Z(4'd2)
	)
	Velocity_Cache_3_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[34*3*DATA_WIDTH-1:33*3*DATA_WIDTH])
	);
	Velocity_Cache_3_1_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd3),
		.CELL_Y(4'd1),
		.CELL_Z(4'd3)
	)
	Velocity_Cache_3_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[35*3*DATA_WIDTH-1:34*3*DATA_WIDTH])
	);
	Velocity_Cache_3_1_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd3),
		.CELL_Y(4'd1),
		.CELL_Z(4'd4)
	)
	Velocity_Cache_3_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[36*3*DATA_WIDTH-1:35*3*DATA_WIDTH])
	);
	Velocity_Cache_3_2_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd3),
		.CELL_Y(4'd2),
		.CELL_Z(4'd1)
	)
	Velocity_Cache_3_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[37*3*DATA_WIDTH-1:36*3*DATA_WIDTH])
	);
	Velocity_Cache_3_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd3),
		.CELL_Y(4'd2),
		.CELL_Z(4'd2)
	)
	Velocity_Cache_3_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[38*3*DATA_WIDTH-1:37*3*DATA_WIDTH])
	);
	Velocity_Cache_3_2_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd3),
		.CELL_Y(4'd2),
		.CELL_Z(4'd3)
	)
	Velocity_Cache_3_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[39*3*DATA_WIDTH-1:38*3*DATA_WIDTH])
	);
	Velocity_Cache_3_2_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd3),
		.CELL_Y(4'd2),
		.CELL_Z(4'd4)
	)
	Velocity_Cache_3_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[40*3*DATA_WIDTH-1:39*3*DATA_WIDTH])
	);
	Velocity_Cache_3_3_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd3),
		.CELL_Y(4'd3),
		.CELL_Z(4'd1)
	)
	Velocity_Cache_3_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[41*3*DATA_WIDTH-1:40*3*DATA_WIDTH])
	);
	Velocity_Cache_3_3_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd3),
		.CELL_Y(4'd3),
		.CELL_Z(4'd2)
	)
	Velocity_Cache_3_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[42*3*DATA_WIDTH-1:41*3*DATA_WIDTH])
	);
	Velocity_Cache_3_3_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd3),
		.CELL_Y(4'd3),
		.CELL_Z(4'd3)
	)
	Velocity_Cache_3_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[43*3*DATA_WIDTH-1:42*3*DATA_WIDTH])
	);
	Velocity_Cache_3_3_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd3),
		.CELL_Y(4'd3),
		.CELL_Z(4'd4)
	)
	Velocity_Cache_3_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[44*3*DATA_WIDTH-1:43*3*DATA_WIDTH])
	);
	Velocity_Cache_3_4_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd3),
		.CELL_Y(4'd4),
		.CELL_Z(4'd1)
	)
	Velocity_Cache_3_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[45*3*DATA_WIDTH-1:44*3*DATA_WIDTH])
	);
	Velocity_Cache_3_4_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd3),
		.CELL_Y(4'd4),
		.CELL_Z(4'd2)
	)
	Velocity_Cache_3_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[46*3*DATA_WIDTH-1:45*3*DATA_WIDTH])
	);
	Velocity_Cache_3_4_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd3),
		.CELL_Y(4'd4),
		.CELL_Z(4'd3)
	)
	Velocity_Cache_3_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[47*3*DATA_WIDTH-1:46*3*DATA_WIDTH])
	);
	Velocity_Cache_3_4_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd3),
		.CELL_Y(4'd4),
		.CELL_Z(4'd4)
	)
	Velocity_Cache_3_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[48*3*DATA_WIDTH-1:47*3*DATA_WIDTH])
	);
	Velocity_Cache_4_1_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd4),
		.CELL_Y(4'd1),
		.CELL_Z(4'd1)
	)
	Velocity_Cache_4_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[49*3*DATA_WIDTH-1:48*3*DATA_WIDTH])
	);
	Velocity_Cache_4_1_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd4),
		.CELL_Y(4'd1),
		.CELL_Z(4'd2)
	)
	Velocity_Cache_4_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[50*3*DATA_WIDTH-1:49*3*DATA_WIDTH])
	);
	Velocity_Cache_4_1_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd4),
		.CELL_Y(4'd1),
		.CELL_Z(4'd3)
	)
	Velocity_Cache_4_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[51*3*DATA_WIDTH-1:50*3*DATA_WIDTH])
	);
	Velocity_Cache_4_1_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd4),
		.CELL_Y(4'd1),
		.CELL_Z(4'd4)
	)
	Velocity_Cache_4_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[52*3*DATA_WIDTH-1:51*3*DATA_WIDTH])
	);
	Velocity_Cache_4_2_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd4),
		.CELL_Y(4'd2),
		.CELL_Z(4'd1)
	)
	Velocity_Cache_4_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[53*3*DATA_WIDTH-1:52*3*DATA_WIDTH])
	);
	Velocity_Cache_4_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd4),
		.CELL_Y(4'd2),
		.CELL_Z(4'd2)
	)
	Velocity_Cache_4_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[54*3*DATA_WIDTH-1:53*3*DATA_WIDTH])
	);
	Velocity_Cache_4_2_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd4),
		.CELL_Y(4'd2),
		.CELL_Z(4'd3)
	)
	Velocity_Cache_4_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[55*3*DATA_WIDTH-1:54*3*DATA_WIDTH])
	);
	Velocity_Cache_4_2_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd4),
		.CELL_Y(4'd2),
		.CELL_Z(4'd4)
	)
	Velocity_Cache_4_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[56*3*DATA_WIDTH-1:55*3*DATA_WIDTH])
	);
	Velocity_Cache_4_3_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd4),
		.CELL_Y(4'd3),
		.CELL_Z(4'd1)
	)
	Velocity_Cache_4_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[57*3*DATA_WIDTH-1:56*3*DATA_WIDTH])
	);
	Velocity_Cache_4_3_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd4),
		.CELL_Y(4'd3),
		.CELL_Z(4'd2)
	)
	Velocity_Cache_4_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[58*3*DATA_WIDTH-1:57*3*DATA_WIDTH])
	);
	Velocity_Cache_4_3_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd4),
		.CELL_Y(4'd3),
		.CELL_Z(4'd3)
	)
	Velocity_Cache_4_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[59*3*DATA_WIDTH-1:58*3*DATA_WIDTH])
	);
	Velocity_Cache_4_3_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd4),
		.CELL_Y(4'd3),
		.CELL_Z(4'd4)
	)
	Velocity_Cache_4_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[60*3*DATA_WIDTH-1:59*3*DATA_WIDTH])
	);
	Velocity_Cache_4_4_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd4),
		.CELL_Y(4'd4),
		.CELL_Z(4'd1)
	)
	Velocity_Cache_4_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[61*3*DATA_WIDTH-1:60*3*DATA_WIDTH])
	);
	Velocity_Cache_4_4_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd4),
		.CELL_Y(4'd4),
		.CELL_Z(4'd2)
	)
	Velocity_Cache_4_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[62*3*DATA_WIDTH-1:61*3*DATA_WIDTH])
	);
	Velocity_Cache_4_4_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd4),
		.CELL_Y(4'd4),
		.CELL_Z(4'd3)
	)
	Velocity_Cache_4_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[63*3*DATA_WIDTH-1:62*3*DATA_WIDTH])
	);
	Velocity_Cache_4_4_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4'd4),
		.CELL_Y(4'd4),
		.CELL_Z(4'd4)
	)
	Velocity_Cache_4_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(Motion_Update_velocity_data[64*3*DATA_WIDTH-1:63*3*DATA_WIDTH])
	);
	
endmodule