/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Module: fp_atan2.v
//
//	Function:
//				Wrapper on top of FP_ATAN, to meet the port configuration in the old design
//
// Dependency:
//				FP_ATAN.v
//
// Latency: 85 cycles
//
//
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module fp_atan2
#(
	parameter DATA_WIDTH = 32
)
(
	input clk,
	input rst,
	input [DATA_WIDTH-1:0] in1,
	input [DATA_WIDTH-1:0] in2,
	output [DATA_WIDTH-1:0] result
);

	FP_ATAN FP_ATAN
	(
		.clk(clk),
		.areset(rst),
		.a(in1),
		.b(in2),
		.q(result)
	);

endmodule
