/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Takes in read addresses of local generators, and map to global cells based on the enable bits.
// If a position cache is read requested by multiple pipelines, the arbiter will resolve the conflict with Round-Robin
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module Local_global_mapping
#(
	parameter NUM_NEIGHBOR_CELLS		= 13,
	parameter NUM_PIPELINES				= 16,
	parameter CELL_ADDR_WIDTH			= 7,
	parameter CELL_ID_WIDTH				= 3,
	parameter NUM_FILTER					= 8,
	parameter TOTAL_CELL_NUM			= 64,
	parameter RDADDR_ARBITER_SIZE		= 5,
	parameter RDADDR_ARBITER_BOTTOM_SIZE = 4,
	parameter RDADDR_ARBITER_MSB		= 16,
	parameter PARTICLE_ID_WIDTH		= CELL_ID_WIDTH*3+CELL_ADDR_WIDTH,
	parameter DATA_WIDTH					= 32
)
(
	input clk,
	input rst,
	input [CELL_ID_WIDTH-1:0] cellz,
	input [NUM_PIPELINES*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:0] Local_FSM_to_Cell_read_addr,
	input [NUM_PIPELINES*(NUM_NEIGHBOR_CELLS+1)-1:0] Local_enable_reading,
	input [TOTAL_CELL_NUM*3*DATA_WIDTH-1:0] Position_Cache_readout_position,
	
	// send to All_Position_Caches
	output [TOTAL_CELL_NUM-1:0] enable_reading,
	output [TOTAL_CELL_NUM*CELL_ADDR_WIDTH-1:0] FSM_to_Cell_read_addr,
	output [NUM_PIPELINES*(NUM_NEIGHBOR_CELLS+1)-1:0] Cell_to_FSM_read_success_bit,
	output [NUM_PIPELINES*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH-1:0] cells_to_pipeline
);
reg [TOTAL_CELL_NUM-1:0] reg_enable_reading;
assign enable_reading = reg_enable_reading;

reg [NUM_PIPELINES*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH-1:0] reg_cells_to_pipeline;
assign cells_to_pipeline = reg_cells_to_pipeline;

always@(*)
	begin
	if (rst)
		begin
		reg_enable_reading = 0;
		reg_cells_to_pipeline = 0;
		end
	else
		begin
		
		// Mapping
		case (cellz)
			1:
				begin
				reg_enable_reading[0] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+0] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+12]);
				reg_enable_reading[1] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+1] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+13]);
				reg_enable_reading[2] <= 0;
				reg_enable_reading[3] <= (Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+2] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+11]);
				reg_enable_reading[4] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+0] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+6]);
				reg_enable_reading[5] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+1] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+7]);
				reg_enable_reading[6] <= 0;
				reg_enable_reading[7] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+2] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+5]);
				reg_enable_reading[8] <= (Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+0] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+6]);
				reg_enable_reading[9] <= (Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+1] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+7]);
				reg_enable_reading[10] <= 0;
				reg_enable_reading[11] <= (Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+2] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+5]);
				reg_enable_reading[12] <= (Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+0] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+9]);
				reg_enable_reading[13] <= (Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+1] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+10]);
				reg_enable_reading[14] <= 0;
				reg_enable_reading[15] <= (Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+2] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+8]);
				reg_enable_reading[16] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+0] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+3]);
				reg_enable_reading[17] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+1] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+4]);
				reg_enable_reading[18] <= 0;
				reg_enable_reading[19] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[20] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[21] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[22] <= 0;
				reg_enable_reading[23] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[24] <= (Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[25] <= (Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[26] <= 0;
				reg_enable_reading[27] <= (Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[28] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[29] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[30] <= 0;
				reg_enable_reading[31] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[32] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+0] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+3]);
				reg_enable_reading[33] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+1] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+4]);
				reg_enable_reading[34] <= 0;
				reg_enable_reading[35] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[36] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[37] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[38] <= 0;
				reg_enable_reading[39] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[40] <= (Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[41] <= (Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[42] <= 0;
				reg_enable_reading[43] <= (Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[44] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[45] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[46] <= 0;
				reg_enable_reading[47] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[48] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+0] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+3]);
				reg_enable_reading[49] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+1] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+4]);
				reg_enable_reading[50] <= 0;
				reg_enable_reading[51] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[52] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[53] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[54] <= 0;
				reg_enable_reading[55] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[56] <= (Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[57] <= (Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[58] <= 0;
				reg_enable_reading[59] <= (Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[60] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[61] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[62] <= 0;
				reg_enable_reading[63] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[12*3*DATA_WIDTH-1:11*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[9*3*DATA_WIDTH-1:8*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[10*3*DATA_WIDTH-1:9*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[28*3*DATA_WIDTH-1:27*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[25*3*DATA_WIDTH-1:24*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[26*3*DATA_WIDTH-1:25*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[9*3*DATA_WIDTH-1:8*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[10*3*DATA_WIDTH-1:9*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[16*3*DATA_WIDTH-1:15*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[13*3*DATA_WIDTH-1:12*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[14*3*DATA_WIDTH-1:13*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[28*3*DATA_WIDTH-1:27*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[25*3*DATA_WIDTH-1:24*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[26*3*DATA_WIDTH-1:25*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[13*3*DATA_WIDTH-1:12*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[14*3*DATA_WIDTH-1:13*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[28*3*DATA_WIDTH-1:27*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[25*3*DATA_WIDTH-1:24*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[26*3*DATA_WIDTH-1:25*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[48*3*DATA_WIDTH-1:47*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[45*3*DATA_WIDTH-1:44*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[46*3*DATA_WIDTH-1:45*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[36*3*DATA_WIDTH-1:35*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[33*3*DATA_WIDTH-1:32*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[34*3*DATA_WIDTH-1:33*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[40*3*DATA_WIDTH-1:39*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[37*3*DATA_WIDTH-1:36*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[38*3*DATA_WIDTH-1:37*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[28*3*DATA_WIDTH-1:27*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[25*3*DATA_WIDTH-1:24*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[26*3*DATA_WIDTH-1:25*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[36*3*DATA_WIDTH-1:35*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[33*3*DATA_WIDTH-1:32*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[34*3*DATA_WIDTH-1:33*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[40*3*DATA_WIDTH-1:39*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[37*3*DATA_WIDTH-1:36*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[38*3*DATA_WIDTH-1:37*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[44*3*DATA_WIDTH-1:43*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[41*3*DATA_WIDTH-1:40*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[42*3*DATA_WIDTH-1:41*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[25*3*DATA_WIDTH-1:24*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[26*3*DATA_WIDTH-1:25*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[40*3*DATA_WIDTH-1:39*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[37*3*DATA_WIDTH-1:36*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[38*3*DATA_WIDTH-1:37*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[44*3*DATA_WIDTH-1:43*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[41*3*DATA_WIDTH-1:40*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[42*3*DATA_WIDTH-1:41*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[48*3*DATA_WIDTH-1:47*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[45*3*DATA_WIDTH-1:44*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[46*3*DATA_WIDTH-1:45*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[44*3*DATA_WIDTH-1:43*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[41*3*DATA_WIDTH-1:40*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[42*3*DATA_WIDTH-1:41*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[48*3*DATA_WIDTH-1:47*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[45*3*DATA_WIDTH-1:44*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[46*3*DATA_WIDTH-1:45*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[36*3*DATA_WIDTH-1:35*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[33*3*DATA_WIDTH-1:32*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[34*3*DATA_WIDTH-1:33*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[33*3*DATA_WIDTH-1:32*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[34*3*DATA_WIDTH-1:33*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[40*3*DATA_WIDTH-1:39*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[37*3*DATA_WIDTH-1:36*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[38*3*DATA_WIDTH-1:37*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[64*3*DATA_WIDTH-1:63*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[61*3*DATA_WIDTH-1:60*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[62*3*DATA_WIDTH-1:61*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[52*3*DATA_WIDTH-1:51*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[49*3*DATA_WIDTH-1:48*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[50*3*DATA_WIDTH-1:49*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[56*3*DATA_WIDTH-1:55*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[53*3*DATA_WIDTH-1:52*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[54*3*DATA_WIDTH-1:53*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[37*3*DATA_WIDTH-1:36*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[38*3*DATA_WIDTH-1:37*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[44*3*DATA_WIDTH-1:43*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[41*3*DATA_WIDTH-1:40*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[42*3*DATA_WIDTH-1:41*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[52*3*DATA_WIDTH-1:51*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[49*3*DATA_WIDTH-1:48*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[50*3*DATA_WIDTH-1:49*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[56*3*DATA_WIDTH-1:55*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[53*3*DATA_WIDTH-1:52*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[54*3*DATA_WIDTH-1:53*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[60*3*DATA_WIDTH-1:59*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[57*3*DATA_WIDTH-1:56*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[58*3*DATA_WIDTH-1:57*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[41*3*DATA_WIDTH-1:40*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[42*3*DATA_WIDTH-1:41*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[48*3*DATA_WIDTH-1:47*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[45*3*DATA_WIDTH-1:44*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[46*3*DATA_WIDTH-1:45*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[56*3*DATA_WIDTH-1:55*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[53*3*DATA_WIDTH-1:52*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[54*3*DATA_WIDTH-1:53*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[60*3*DATA_WIDTH-1:59*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[57*3*DATA_WIDTH-1:56*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[58*3*DATA_WIDTH-1:57*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[64*3*DATA_WIDTH-1:63*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[61*3*DATA_WIDTH-1:60*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[62*3*DATA_WIDTH-1:61*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[45*3*DATA_WIDTH-1:44*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[46*3*DATA_WIDTH-1:45*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[36*3*DATA_WIDTH-1:35*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[33*3*DATA_WIDTH-1:32*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[34*3*DATA_WIDTH-1:33*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[60*3*DATA_WIDTH-1:59*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[57*3*DATA_WIDTH-1:56*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[58*3*DATA_WIDTH-1:57*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[64*3*DATA_WIDTH-1:63*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[61*3*DATA_WIDTH-1:60*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[62*3*DATA_WIDTH-1:61*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[52*3*DATA_WIDTH-1:51*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[49*3*DATA_WIDTH-1:48*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[50*3*DATA_WIDTH-1:49*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[49*3*DATA_WIDTH-1:48*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[50*3*DATA_WIDTH-1:49*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[56*3*DATA_WIDTH-1:55*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[53*3*DATA_WIDTH-1:52*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[54*3*DATA_WIDTH-1:53*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[16*3*DATA_WIDTH-1:15*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[13*3*DATA_WIDTH-1:12*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[14*3*DATA_WIDTH-1:13*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[53*3*DATA_WIDTH-1:52*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[54*3*DATA_WIDTH-1:53*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[60*3*DATA_WIDTH-1:59*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[57*3*DATA_WIDTH-1:56*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[58*3*DATA_WIDTH-1:57*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[12*3*DATA_WIDTH-1:11*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[9*3*DATA_WIDTH-1:8*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[10*3*DATA_WIDTH-1:9*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[57*3*DATA_WIDTH-1:56*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[58*3*DATA_WIDTH-1:57*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[64*3*DATA_WIDTH-1:63*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[61*3*DATA_WIDTH-1:60*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[62*3*DATA_WIDTH-1:61*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[12*3*DATA_WIDTH-1:11*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[9*3*DATA_WIDTH-1:8*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[10*3*DATA_WIDTH-1:9*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[16*3*DATA_WIDTH-1:15*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[13*3*DATA_WIDTH-1:12*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[14*3*DATA_WIDTH-1:13*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[61*3*DATA_WIDTH-1:60*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[62*3*DATA_WIDTH-1:61*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[52*3*DATA_WIDTH-1:51*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[49*3*DATA_WIDTH-1:48*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[50*3*DATA_WIDTH-1:49*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[12*3*DATA_WIDTH-1:11*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[9*3*DATA_WIDTH-1:8*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[10*3*DATA_WIDTH-1:9*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[16*3*DATA_WIDTH-1:15*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[13*3*DATA_WIDTH-1:12*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[14*3*DATA_WIDTH-1:13*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH];
				end
			2:
				begin
				reg_enable_reading[0] <= (Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+2] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+11]);
				reg_enable_reading[1] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+0] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+12]);
				reg_enable_reading[2] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+1] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+13]);
				reg_enable_reading[3] <= 0;
				reg_enable_reading[4] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+2] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+5]);
				reg_enable_reading[5] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+0] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+6]);
				reg_enable_reading[6] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+1] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+7]);
				reg_enable_reading[7] <= 0;
				reg_enable_reading[8] <= (Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+2] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+5]);
				reg_enable_reading[9] <= (Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+0] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+6]);
				reg_enable_reading[10] <= (Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+1] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+7]);
				reg_enable_reading[11] <= 0;
				reg_enable_reading[12] <= (Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+2] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+8]);
				reg_enable_reading[13] <= (Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+0] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+9]);
				reg_enable_reading[14] <= (Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+1] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+10]);
				reg_enable_reading[15] <= 0;
				reg_enable_reading[16] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[17] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+0] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+3]);
				reg_enable_reading[18] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+1] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+4]);
				reg_enable_reading[19] <= 0;
				reg_enable_reading[20] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[21] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[22] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[23] <= 0;
				reg_enable_reading[24] <= (Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[25] <= (Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[26] <= (Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[27] <= 0;
				reg_enable_reading[28] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[29] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[30] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[31] <= 0;
				reg_enable_reading[32] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[33] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+0] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+3]);
				reg_enable_reading[34] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+1] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+4]);
				reg_enable_reading[35] <= 0;
				reg_enable_reading[36] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[37] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[38] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[39] <= 0;
				reg_enable_reading[40] <= (Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[41] <= (Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[42] <= (Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[43] <= 0;
				reg_enable_reading[44] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[45] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[46] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[47] <= 0;
				reg_enable_reading[48] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[49] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+0] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+3]);
				reg_enable_reading[50] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+1] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+4]);
				reg_enable_reading[51] <= 0;
				reg_enable_reading[52] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[53] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[54] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[55] <= 0;
				reg_enable_reading[56] <= (Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[57] <= (Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[58] <= (Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[59] <= 0;
				reg_enable_reading[60] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[61] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[62] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[63] <= 0;
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[9*3*DATA_WIDTH-1:8*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[10*3*DATA_WIDTH-1:9*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[11*3*DATA_WIDTH-1:10*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[25*3*DATA_WIDTH-1:24*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[26*3*DATA_WIDTH-1:25*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[27*3*DATA_WIDTH-1:26*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[10*3*DATA_WIDTH-1:9*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[11*3*DATA_WIDTH-1:10*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[13*3*DATA_WIDTH-1:12*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[14*3*DATA_WIDTH-1:13*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[15*3*DATA_WIDTH-1:14*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[25*3*DATA_WIDTH-1:24*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[26*3*DATA_WIDTH-1:25*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[27*3*DATA_WIDTH-1:26*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[14*3*DATA_WIDTH-1:13*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[15*3*DATA_WIDTH-1:14*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[25*3*DATA_WIDTH-1:24*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[26*3*DATA_WIDTH-1:25*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[27*3*DATA_WIDTH-1:26*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[45*3*DATA_WIDTH-1:44*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[46*3*DATA_WIDTH-1:45*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[47*3*DATA_WIDTH-1:46*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[33*3*DATA_WIDTH-1:32*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[34*3*DATA_WIDTH-1:33*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[35*3*DATA_WIDTH-1:34*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[37*3*DATA_WIDTH-1:36*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[38*3*DATA_WIDTH-1:37*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[39*3*DATA_WIDTH-1:38*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[25*3*DATA_WIDTH-1:24*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[26*3*DATA_WIDTH-1:25*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[27*3*DATA_WIDTH-1:26*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[33*3*DATA_WIDTH-1:32*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[34*3*DATA_WIDTH-1:33*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[35*3*DATA_WIDTH-1:34*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[37*3*DATA_WIDTH-1:36*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[38*3*DATA_WIDTH-1:37*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[39*3*DATA_WIDTH-1:38*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[41*3*DATA_WIDTH-1:40*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[42*3*DATA_WIDTH-1:41*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[43*3*DATA_WIDTH-1:42*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[26*3*DATA_WIDTH-1:25*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[27*3*DATA_WIDTH-1:26*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[37*3*DATA_WIDTH-1:36*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[38*3*DATA_WIDTH-1:37*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[39*3*DATA_WIDTH-1:38*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[41*3*DATA_WIDTH-1:40*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[42*3*DATA_WIDTH-1:41*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[43*3*DATA_WIDTH-1:42*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[45*3*DATA_WIDTH-1:44*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[46*3*DATA_WIDTH-1:45*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[47*3*DATA_WIDTH-1:46*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[41*3*DATA_WIDTH-1:40*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[42*3*DATA_WIDTH-1:41*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[43*3*DATA_WIDTH-1:42*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[45*3*DATA_WIDTH-1:44*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[46*3*DATA_WIDTH-1:45*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[47*3*DATA_WIDTH-1:46*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[33*3*DATA_WIDTH-1:32*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[34*3*DATA_WIDTH-1:33*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[35*3*DATA_WIDTH-1:34*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[34*3*DATA_WIDTH-1:33*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[35*3*DATA_WIDTH-1:34*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[37*3*DATA_WIDTH-1:36*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[38*3*DATA_WIDTH-1:37*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[39*3*DATA_WIDTH-1:38*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[61*3*DATA_WIDTH-1:60*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[62*3*DATA_WIDTH-1:61*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[63*3*DATA_WIDTH-1:62*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[49*3*DATA_WIDTH-1:48*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[50*3*DATA_WIDTH-1:49*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[51*3*DATA_WIDTH-1:50*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[53*3*DATA_WIDTH-1:52*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[54*3*DATA_WIDTH-1:53*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[55*3*DATA_WIDTH-1:54*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[38*3*DATA_WIDTH-1:37*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[39*3*DATA_WIDTH-1:38*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[41*3*DATA_WIDTH-1:40*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[42*3*DATA_WIDTH-1:41*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[43*3*DATA_WIDTH-1:42*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[49*3*DATA_WIDTH-1:48*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[50*3*DATA_WIDTH-1:49*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[51*3*DATA_WIDTH-1:50*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[53*3*DATA_WIDTH-1:52*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[54*3*DATA_WIDTH-1:53*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[55*3*DATA_WIDTH-1:54*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[57*3*DATA_WIDTH-1:56*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[58*3*DATA_WIDTH-1:57*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[59*3*DATA_WIDTH-1:58*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[42*3*DATA_WIDTH-1:41*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[43*3*DATA_WIDTH-1:42*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[45*3*DATA_WIDTH-1:44*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[46*3*DATA_WIDTH-1:45*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[47*3*DATA_WIDTH-1:46*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[53*3*DATA_WIDTH-1:52*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[54*3*DATA_WIDTH-1:53*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[55*3*DATA_WIDTH-1:54*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[57*3*DATA_WIDTH-1:56*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[58*3*DATA_WIDTH-1:57*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[59*3*DATA_WIDTH-1:58*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[61*3*DATA_WIDTH-1:60*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[62*3*DATA_WIDTH-1:61*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[63*3*DATA_WIDTH-1:62*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[46*3*DATA_WIDTH-1:45*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[47*3*DATA_WIDTH-1:46*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[33*3*DATA_WIDTH-1:32*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[34*3*DATA_WIDTH-1:33*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[35*3*DATA_WIDTH-1:34*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[57*3*DATA_WIDTH-1:56*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[58*3*DATA_WIDTH-1:57*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[59*3*DATA_WIDTH-1:58*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[61*3*DATA_WIDTH-1:60*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[62*3*DATA_WIDTH-1:61*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[63*3*DATA_WIDTH-1:62*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[49*3*DATA_WIDTH-1:48*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[50*3*DATA_WIDTH-1:49*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[51*3*DATA_WIDTH-1:50*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[50*3*DATA_WIDTH-1:49*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[51*3*DATA_WIDTH-1:50*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[53*3*DATA_WIDTH-1:52*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[54*3*DATA_WIDTH-1:53*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[55*3*DATA_WIDTH-1:54*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[13*3*DATA_WIDTH-1:12*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[14*3*DATA_WIDTH-1:13*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[15*3*DATA_WIDTH-1:14*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[54*3*DATA_WIDTH-1:53*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[55*3*DATA_WIDTH-1:54*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[57*3*DATA_WIDTH-1:56*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[58*3*DATA_WIDTH-1:57*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[59*3*DATA_WIDTH-1:58*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[9*3*DATA_WIDTH-1:8*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[10*3*DATA_WIDTH-1:9*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[11*3*DATA_WIDTH-1:10*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[58*3*DATA_WIDTH-1:57*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[59*3*DATA_WIDTH-1:58*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[61*3*DATA_WIDTH-1:60*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[62*3*DATA_WIDTH-1:61*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[63*3*DATA_WIDTH-1:62*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[9*3*DATA_WIDTH-1:8*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[10*3*DATA_WIDTH-1:9*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[11*3*DATA_WIDTH-1:10*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[13*3*DATA_WIDTH-1:12*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[14*3*DATA_WIDTH-1:13*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[15*3*DATA_WIDTH-1:14*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[62*3*DATA_WIDTH-1:61*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[63*3*DATA_WIDTH-1:62*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[49*3*DATA_WIDTH-1:48*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[50*3*DATA_WIDTH-1:49*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[51*3*DATA_WIDTH-1:50*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[9*3*DATA_WIDTH-1:8*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[10*3*DATA_WIDTH-1:9*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[11*3*DATA_WIDTH-1:10*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[13*3*DATA_WIDTH-1:12*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[14*3*DATA_WIDTH-1:13*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[15*3*DATA_WIDTH-1:14*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH];
				end
			3:
				begin
				reg_enable_reading[0] <= 0;
				reg_enable_reading[1] <= (Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+2] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+11]);
				reg_enable_reading[2] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+0] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+12]);
				reg_enable_reading[3] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+1] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+13]);
				reg_enable_reading[4] <= 0;
				reg_enable_reading[5] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+2] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+5]);
				reg_enable_reading[6] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+0] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+6]);
				reg_enable_reading[7] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+1] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+7]);
				reg_enable_reading[8] <= 0;
				reg_enable_reading[9] <= (Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+2] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+5]);
				reg_enable_reading[10] <= (Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+0] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+6]);
				reg_enable_reading[11] <= (Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+1] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+7]);
				reg_enable_reading[12] <= 0;
				reg_enable_reading[13] <= (Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+2] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+8]);
				reg_enable_reading[14] <= (Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+0] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+9]);
				reg_enable_reading[15] <= (Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+1] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+10]);
				reg_enable_reading[16] <= 0;
				reg_enable_reading[17] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[18] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+0] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+3]);
				reg_enable_reading[19] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+1] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+4]);
				reg_enable_reading[20] <= 0;
				reg_enable_reading[21] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[22] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[23] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[24] <= 0;
				reg_enable_reading[25] <= (Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[26] <= (Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[27] <= (Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[28] <= 0;
				reg_enable_reading[29] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[30] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[31] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[32] <= 0;
				reg_enable_reading[33] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[34] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+0] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+3]);
				reg_enable_reading[35] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+1] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+4]);
				reg_enable_reading[36] <= 0;
				reg_enable_reading[37] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[38] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[39] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[40] <= 0;
				reg_enable_reading[41] <= (Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[42] <= (Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[43] <= (Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[44] <= 0;
				reg_enable_reading[45] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[46] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[47] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[48] <= 0;
				reg_enable_reading[49] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[50] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+0] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+3]);
				reg_enable_reading[51] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+1] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+4]);
				reg_enable_reading[52] <= 0;
				reg_enable_reading[53] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[54] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[55] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[56] <= 0;
				reg_enable_reading[57] <= (Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[58] <= (Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[59] <= (Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[60] <= 0;
				reg_enable_reading[61] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[62] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[63] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[10*3*DATA_WIDTH-1:9*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[11*3*DATA_WIDTH-1:10*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[12*3*DATA_WIDTH-1:11*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[26*3*DATA_WIDTH-1:25*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[27*3*DATA_WIDTH-1:26*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[28*3*DATA_WIDTH-1:27*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[11*3*DATA_WIDTH-1:10*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[12*3*DATA_WIDTH-1:11*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[14*3*DATA_WIDTH-1:13*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[15*3*DATA_WIDTH-1:14*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[16*3*DATA_WIDTH-1:15*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[26*3*DATA_WIDTH-1:25*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[27*3*DATA_WIDTH-1:26*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[28*3*DATA_WIDTH-1:27*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[15*3*DATA_WIDTH-1:14*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[16*3*DATA_WIDTH-1:15*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[26*3*DATA_WIDTH-1:25*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[27*3*DATA_WIDTH-1:26*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[28*3*DATA_WIDTH-1:27*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[46*3*DATA_WIDTH-1:45*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[47*3*DATA_WIDTH-1:46*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[48*3*DATA_WIDTH-1:47*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[34*3*DATA_WIDTH-1:33*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[35*3*DATA_WIDTH-1:34*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[36*3*DATA_WIDTH-1:35*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[38*3*DATA_WIDTH-1:37*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[39*3*DATA_WIDTH-1:38*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[40*3*DATA_WIDTH-1:39*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[26*3*DATA_WIDTH-1:25*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[27*3*DATA_WIDTH-1:26*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[28*3*DATA_WIDTH-1:27*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[34*3*DATA_WIDTH-1:33*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[35*3*DATA_WIDTH-1:34*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[36*3*DATA_WIDTH-1:35*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[38*3*DATA_WIDTH-1:37*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[39*3*DATA_WIDTH-1:38*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[40*3*DATA_WIDTH-1:39*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[42*3*DATA_WIDTH-1:41*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[43*3*DATA_WIDTH-1:42*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[44*3*DATA_WIDTH-1:43*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[27*3*DATA_WIDTH-1:26*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[28*3*DATA_WIDTH-1:27*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[38*3*DATA_WIDTH-1:37*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[39*3*DATA_WIDTH-1:38*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[40*3*DATA_WIDTH-1:39*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[42*3*DATA_WIDTH-1:41*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[43*3*DATA_WIDTH-1:42*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[44*3*DATA_WIDTH-1:43*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[46*3*DATA_WIDTH-1:45*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[47*3*DATA_WIDTH-1:46*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[48*3*DATA_WIDTH-1:47*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[42*3*DATA_WIDTH-1:41*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[43*3*DATA_WIDTH-1:42*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[44*3*DATA_WIDTH-1:43*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[46*3*DATA_WIDTH-1:45*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[47*3*DATA_WIDTH-1:46*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[48*3*DATA_WIDTH-1:47*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[34*3*DATA_WIDTH-1:33*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[35*3*DATA_WIDTH-1:34*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[36*3*DATA_WIDTH-1:35*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[35*3*DATA_WIDTH-1:34*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[36*3*DATA_WIDTH-1:35*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[38*3*DATA_WIDTH-1:37*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[39*3*DATA_WIDTH-1:38*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[40*3*DATA_WIDTH-1:39*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[62*3*DATA_WIDTH-1:61*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[63*3*DATA_WIDTH-1:62*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[64*3*DATA_WIDTH-1:63*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[50*3*DATA_WIDTH-1:49*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[51*3*DATA_WIDTH-1:50*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[52*3*DATA_WIDTH-1:51*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[54*3*DATA_WIDTH-1:53*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[55*3*DATA_WIDTH-1:54*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[56*3*DATA_WIDTH-1:55*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[39*3*DATA_WIDTH-1:38*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[40*3*DATA_WIDTH-1:39*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[42*3*DATA_WIDTH-1:41*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[43*3*DATA_WIDTH-1:42*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[44*3*DATA_WIDTH-1:43*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[50*3*DATA_WIDTH-1:49*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[51*3*DATA_WIDTH-1:50*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[52*3*DATA_WIDTH-1:51*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[54*3*DATA_WIDTH-1:53*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[55*3*DATA_WIDTH-1:54*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[56*3*DATA_WIDTH-1:55*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[58*3*DATA_WIDTH-1:57*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[59*3*DATA_WIDTH-1:58*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[60*3*DATA_WIDTH-1:59*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[43*3*DATA_WIDTH-1:42*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[44*3*DATA_WIDTH-1:43*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[46*3*DATA_WIDTH-1:45*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[47*3*DATA_WIDTH-1:46*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[48*3*DATA_WIDTH-1:47*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[54*3*DATA_WIDTH-1:53*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[55*3*DATA_WIDTH-1:54*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[56*3*DATA_WIDTH-1:55*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[58*3*DATA_WIDTH-1:57*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[59*3*DATA_WIDTH-1:58*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[60*3*DATA_WIDTH-1:59*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[62*3*DATA_WIDTH-1:61*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[63*3*DATA_WIDTH-1:62*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[64*3*DATA_WIDTH-1:63*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[47*3*DATA_WIDTH-1:46*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[48*3*DATA_WIDTH-1:47*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[34*3*DATA_WIDTH-1:33*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[35*3*DATA_WIDTH-1:34*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[36*3*DATA_WIDTH-1:35*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[58*3*DATA_WIDTH-1:57*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[59*3*DATA_WIDTH-1:58*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[60*3*DATA_WIDTH-1:59*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[62*3*DATA_WIDTH-1:61*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[63*3*DATA_WIDTH-1:62*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[64*3*DATA_WIDTH-1:63*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[50*3*DATA_WIDTH-1:49*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[51*3*DATA_WIDTH-1:50*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[52*3*DATA_WIDTH-1:51*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[51*3*DATA_WIDTH-1:50*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[52*3*DATA_WIDTH-1:51*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[54*3*DATA_WIDTH-1:53*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[55*3*DATA_WIDTH-1:54*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[56*3*DATA_WIDTH-1:55*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[14*3*DATA_WIDTH-1:13*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[15*3*DATA_WIDTH-1:14*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[16*3*DATA_WIDTH-1:15*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[55*3*DATA_WIDTH-1:54*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[56*3*DATA_WIDTH-1:55*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[58*3*DATA_WIDTH-1:57*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[59*3*DATA_WIDTH-1:58*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[60*3*DATA_WIDTH-1:59*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[10*3*DATA_WIDTH-1:9*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[11*3*DATA_WIDTH-1:10*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[12*3*DATA_WIDTH-1:11*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[59*3*DATA_WIDTH-1:58*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[60*3*DATA_WIDTH-1:59*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[62*3*DATA_WIDTH-1:61*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[63*3*DATA_WIDTH-1:62*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[64*3*DATA_WIDTH-1:63*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[10*3*DATA_WIDTH-1:9*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[11*3*DATA_WIDTH-1:10*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[12*3*DATA_WIDTH-1:11*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[14*3*DATA_WIDTH-1:13*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[15*3*DATA_WIDTH-1:14*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[16*3*DATA_WIDTH-1:15*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[63*3*DATA_WIDTH-1:62*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[64*3*DATA_WIDTH-1:63*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[50*3*DATA_WIDTH-1:49*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[51*3*DATA_WIDTH-1:50*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[52*3*DATA_WIDTH-1:51*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[10*3*DATA_WIDTH-1:9*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[11*3*DATA_WIDTH-1:10*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[12*3*DATA_WIDTH-1:11*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[14*3*DATA_WIDTH-1:13*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[15*3*DATA_WIDTH-1:14*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[16*3*DATA_WIDTH-1:15*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH];
				end
			4:
				begin
				reg_enable_reading[0] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+1] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+13]);
				reg_enable_reading[1] <= 0;
				reg_enable_reading[2] <= (Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+2] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+11]);
				reg_enable_reading[3] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+0] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+12]);
				reg_enable_reading[4] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+1] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+7]);
				reg_enable_reading[5] <= 0;
				reg_enable_reading[6] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+2] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+5]);
				reg_enable_reading[7] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+0] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+6]);
				reg_enable_reading[8] <= (Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+1] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+7]);
				reg_enable_reading[9] <= 0;
				reg_enable_reading[10] <= (Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+2] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+5]);
				reg_enable_reading[11] <= (Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+0] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+6]);
				reg_enable_reading[12] <= (Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+1] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+10]);
				reg_enable_reading[13] <= 0;
				reg_enable_reading[14] <= (Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+2] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+8]);
				reg_enable_reading[15] <= (Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+0] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+9]);
				reg_enable_reading[16] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+1] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+4]);
				reg_enable_reading[17] <= 0;
				reg_enable_reading[18] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[19] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+0] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+3]);
				reg_enable_reading[20] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[21] <= 0;
				reg_enable_reading[22] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[23] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[24] <= (Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[25] <= 0;
				reg_enable_reading[26] <= (Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[27] <= (Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[28] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[29] <= 0;
				reg_enable_reading[30] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[31] <= (Local_enable_reading[0*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[32] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+1] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+4]);
				reg_enable_reading[33] <= 0;
				reg_enable_reading[34] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[35] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+0] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+3]);
				reg_enable_reading[36] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[37] <= 0;
				reg_enable_reading[38] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[39] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[40] <= (Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[41] <= 0;
				reg_enable_reading[42] <= (Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[43] <= (Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[44] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[45] <= 0;
				reg_enable_reading[46] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[47] <= (Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[48] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+1] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+4]);
				reg_enable_reading[49] <= 0;
				reg_enable_reading[50] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[51] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+0] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+3]);
				reg_enable_reading[52] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[53] <= 0;
				reg_enable_reading[54] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[55] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[56] <= (Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[57] <= 0;
				reg_enable_reading[58] <= (Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[59] <= (Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_enable_reading[60] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+7] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+13] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+10] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+4] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+1]);
				reg_enable_reading[61] <= 0;
				reg_enable_reading[62] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+5] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+11] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+8] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+2]);
				reg_enable_reading[63] <= (Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)+6] || Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)+12] || Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)+9] || Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)+3] || Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)+0]);
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH];
				reg_cells_to_pipeline[0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[11*3*DATA_WIDTH-1:10*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[12*3*DATA_WIDTH-1:11*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[9*3*DATA_WIDTH-1:8*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[27*3*DATA_WIDTH-1:26*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[28*3*DATA_WIDTH-1:27*3*DATA_WIDTH];
				reg_cells_to_pipeline[1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[25*3*DATA_WIDTH-1:24*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[12*3*DATA_WIDTH-1:11*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[9*3*DATA_WIDTH-1:8*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[15*3*DATA_WIDTH-1:14*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[16*3*DATA_WIDTH-1:15*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[13*3*DATA_WIDTH-1:12*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[27*3*DATA_WIDTH-1:26*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[28*3*DATA_WIDTH-1:27*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[25*3*DATA_WIDTH-1:24*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH];
				reg_cells_to_pipeline[2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[16*3*DATA_WIDTH-1:15*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[13*3*DATA_WIDTH-1:12*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[27*3*DATA_WIDTH-1:26*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[28*3*DATA_WIDTH-1:27*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[25*3*DATA_WIDTH-1:24*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH];
				reg_cells_to_pipeline[3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[47*3*DATA_WIDTH-1:46*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[48*3*DATA_WIDTH-1:47*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[45*3*DATA_WIDTH-1:44*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[35*3*DATA_WIDTH-1:34*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[36*3*DATA_WIDTH-1:35*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[33*3*DATA_WIDTH-1:32*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[39*3*DATA_WIDTH-1:38*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[40*3*DATA_WIDTH-1:39*3*DATA_WIDTH];
				reg_cells_to_pipeline[4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[37*3*DATA_WIDTH-1:36*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[27*3*DATA_WIDTH-1:26*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[28*3*DATA_WIDTH-1:27*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[25*3*DATA_WIDTH-1:24*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[35*3*DATA_WIDTH-1:34*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[36*3*DATA_WIDTH-1:35*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[33*3*DATA_WIDTH-1:32*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[39*3*DATA_WIDTH-1:38*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[40*3*DATA_WIDTH-1:39*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[37*3*DATA_WIDTH-1:36*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[43*3*DATA_WIDTH-1:42*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[44*3*DATA_WIDTH-1:43*3*DATA_WIDTH];
				reg_cells_to_pipeline[5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[41*3*DATA_WIDTH-1:40*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[28*3*DATA_WIDTH-1:27*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[25*3*DATA_WIDTH-1:24*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[39*3*DATA_WIDTH-1:38*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[40*3*DATA_WIDTH-1:39*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[37*3*DATA_WIDTH-1:36*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[43*3*DATA_WIDTH-1:42*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[44*3*DATA_WIDTH-1:43*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[41*3*DATA_WIDTH-1:40*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[47*3*DATA_WIDTH-1:46*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[48*3*DATA_WIDTH-1:47*3*DATA_WIDTH];
				reg_cells_to_pipeline[6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[45*3*DATA_WIDTH-1:44*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[43*3*DATA_WIDTH-1:42*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[44*3*DATA_WIDTH-1:43*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[41*3*DATA_WIDTH-1:40*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[47*3*DATA_WIDTH-1:46*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[48*3*DATA_WIDTH-1:47*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[45*3*DATA_WIDTH-1:44*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[35*3*DATA_WIDTH-1:34*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[36*3*DATA_WIDTH-1:35*3*DATA_WIDTH];
				reg_cells_to_pipeline[7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[33*3*DATA_WIDTH-1:32*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[36*3*DATA_WIDTH-1:35*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[33*3*DATA_WIDTH-1:32*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[39*3*DATA_WIDTH-1:38*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[40*3*DATA_WIDTH-1:39*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[37*3*DATA_WIDTH-1:36*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[63*3*DATA_WIDTH-1:62*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[64*3*DATA_WIDTH-1:63*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[61*3*DATA_WIDTH-1:60*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[51*3*DATA_WIDTH-1:50*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[52*3*DATA_WIDTH-1:51*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[49*3*DATA_WIDTH-1:48*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[55*3*DATA_WIDTH-1:54*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[56*3*DATA_WIDTH-1:55*3*DATA_WIDTH];
				reg_cells_to_pipeline[8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[53*3*DATA_WIDTH-1:52*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[40*3*DATA_WIDTH-1:39*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[37*3*DATA_WIDTH-1:36*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[43*3*DATA_WIDTH-1:42*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[44*3*DATA_WIDTH-1:43*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[41*3*DATA_WIDTH-1:40*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[51*3*DATA_WIDTH-1:50*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[52*3*DATA_WIDTH-1:51*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[49*3*DATA_WIDTH-1:48*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[55*3*DATA_WIDTH-1:54*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[56*3*DATA_WIDTH-1:55*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[53*3*DATA_WIDTH-1:52*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[59*3*DATA_WIDTH-1:58*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[60*3*DATA_WIDTH-1:59*3*DATA_WIDTH];
				reg_cells_to_pipeline[9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[57*3*DATA_WIDTH-1:56*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[44*3*DATA_WIDTH-1:43*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[41*3*DATA_WIDTH-1:40*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[47*3*DATA_WIDTH-1:46*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[48*3*DATA_WIDTH-1:47*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[45*3*DATA_WIDTH-1:44*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[55*3*DATA_WIDTH-1:54*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[56*3*DATA_WIDTH-1:55*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[53*3*DATA_WIDTH-1:52*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[59*3*DATA_WIDTH-1:58*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[60*3*DATA_WIDTH-1:59*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[57*3*DATA_WIDTH-1:56*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[63*3*DATA_WIDTH-1:62*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[64*3*DATA_WIDTH-1:63*3*DATA_WIDTH];
				reg_cells_to_pipeline[10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[61*3*DATA_WIDTH-1:60*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[48*3*DATA_WIDTH-1:47*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[45*3*DATA_WIDTH-1:44*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[35*3*DATA_WIDTH-1:34*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[36*3*DATA_WIDTH-1:35*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[33*3*DATA_WIDTH-1:32*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[59*3*DATA_WIDTH-1:58*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[60*3*DATA_WIDTH-1:59*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[57*3*DATA_WIDTH-1:56*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[63*3*DATA_WIDTH-1:62*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[64*3*DATA_WIDTH-1:63*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[61*3*DATA_WIDTH-1:60*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[51*3*DATA_WIDTH-1:50*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[52*3*DATA_WIDTH-1:51*3*DATA_WIDTH];
				reg_cells_to_pipeline[11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[49*3*DATA_WIDTH-1:48*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[52*3*DATA_WIDTH-1:51*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[49*3*DATA_WIDTH-1:48*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[55*3*DATA_WIDTH-1:54*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[56*3*DATA_WIDTH-1:55*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[53*3*DATA_WIDTH-1:52*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[15*3*DATA_WIDTH-1:14*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[16*3*DATA_WIDTH-1:15*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[13*3*DATA_WIDTH-1:12*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH];
				reg_cells_to_pipeline[12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[56*3*DATA_WIDTH-1:55*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[53*3*DATA_WIDTH-1:52*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[59*3*DATA_WIDTH-1:58*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[60*3*DATA_WIDTH-1:59*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[57*3*DATA_WIDTH-1:56*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[11*3*DATA_WIDTH-1:10*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[12*3*DATA_WIDTH-1:11*3*DATA_WIDTH];
				reg_cells_to_pipeline[13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[9*3*DATA_WIDTH-1:8*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[60*3*DATA_WIDTH-1:59*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[57*3*DATA_WIDTH-1:56*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[63*3*DATA_WIDTH-1:62*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[64*3*DATA_WIDTH-1:63*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[61*3*DATA_WIDTH-1:60*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[11*3*DATA_WIDTH-1:10*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[12*3*DATA_WIDTH-1:11*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[9*3*DATA_WIDTH-1:8*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[15*3*DATA_WIDTH-1:14*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[16*3*DATA_WIDTH-1:15*3*DATA_WIDTH];
				reg_cells_to_pipeline[14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[13*3*DATA_WIDTH-1:12*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+0*3*DATA_WIDTH] <= Position_Cache_readout_position[64*3*DATA_WIDTH-1:63*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+1*3*DATA_WIDTH] <= Position_Cache_readout_position[61*3*DATA_WIDTH-1:60*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+2*3*DATA_WIDTH] <= Position_Cache_readout_position[51*3*DATA_WIDTH-1:50*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+3*3*DATA_WIDTH] <= Position_Cache_readout_position[52*3*DATA_WIDTH-1:51*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+4*3*DATA_WIDTH] <= Position_Cache_readout_position[49*3*DATA_WIDTH-1:48*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+5*3*DATA_WIDTH] <= Position_Cache_readout_position[11*3*DATA_WIDTH-1:10*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+6*3*DATA_WIDTH] <= Position_Cache_readout_position[12*3*DATA_WIDTH-1:11*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+7*3*DATA_WIDTH] <= Position_Cache_readout_position[9*3*DATA_WIDTH-1:8*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+8*3*DATA_WIDTH] <= Position_Cache_readout_position[15*3*DATA_WIDTH-1:14*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+9*3*DATA_WIDTH] <= Position_Cache_readout_position[16*3*DATA_WIDTH-1:15*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+10*3*DATA_WIDTH] <= Position_Cache_readout_position[13*3*DATA_WIDTH-1:12*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+11*3*DATA_WIDTH] <= Position_Cache_readout_position[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+12*3*DATA_WIDTH] <= Position_Cache_readout_position[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH];
				reg_cells_to_pipeline[15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+14*3*DATA_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH+13*3*DATA_WIDTH] <= Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH];
				end
			default:
				begin
				reg_enable_reading = 0;
				reg_cells_to_pipeline = 0;
				end
		endcase
		end
	end
	
Arbitration_Unit
#(
	.NUM_PIPELINES(NUM_PIPELINES),
	.NUM_NEIGHBOR_CELLS(NUM_NEIGHBOR_CELLS),
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.CELL_ID_WIDTH(CELL_ID_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_BOTTOM_SIZE(RDADDR_ARBITER_BOTTOM_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB),
	.TOTAL_CELL_NUM(TOTAL_CELL_NUM)
)
Arbitration_Unit
(
	.clk(clk),
	.rst(rst),
	.cellz(cellz),
	.Local_FSM_to_Cell_read_addr(Local_FSM_to_Cell_read_addr),
	.Local_enable_reading(Local_enable_reading),
	
	.Cell_to_FSM_read_success_bit(Cell_to_FSM_read_success_bit),
	.FSM_to_Cell_read_addr(FSM_to_Cell_read_addr)
);

endmodule