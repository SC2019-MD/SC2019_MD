module Force_Writeback_Arbitration_Unit
#(
	parameter BINARY_222							= 9'b010010010,			// xyz
	parameter BINARY_223							= 9'b010010011,
	parameter BINARY_231							= 9'b010011001,
	parameter BINARY_232							= 9'b010011010,
	parameter BINARY_233							= 9'b010011011,
	parameter BINARY_311							= 9'b011001001,
	parameter BINARY_312							= 9'b011001010,
	parameter BINARY_313							= 9'b011001011,
	parameter BINARY_321							= 9'b011010001,
	parameter BINARY_322							= 9'b011010010,
	parameter BINARY_323							= 9'b011010011,
	parameter BINARY_331							= 9'b011011001,
	parameter BINARY_332							= 9'b011011010,
	parameter BINARY_333							= 9'b011011011,
	parameter NUM_PIPELINES						= 16,
	parameter DATA_WIDTH							= 32,
	parameter CELL_ID_WIDTH						= 3,
	parameter CELL_ADDR_WIDTH					= 7,
	parameter TOTAL_CELL_NUM					= 64,
	parameter PARTICLE_ID_WIDTH				= CELL_ID_WIDTH*3+CELL_ADDR_WIDTH,
	parameter FORCE_WTADDR_ARBITER_SIZE		= 6,
	parameter FORCE_WTADDR_ARBITER_MSB		= 32,
	parameter FORCE_EVAL_FIFO_DATA_WIDTH	= 113,
	parameter FORCE_EVAL_FIFO_DEPTH			= 128,
	parameter FORCE_EVAL_FIFO_ADDR_WIDTH	= 7
)
(
	input clk,
	input rst,
	input [NUM_PIPELINES*FORCE_EVAL_FIFO_DATA_WIDTH-1:0] ref_force_data_from_FIFO,
	input [NUM_PIPELINES*FORCE_EVAL_FIFO_DATA_WIDTH-1:0] neighbor_force_data_from_FIFO_1,
	input [NUM_PIPELINES*FORCE_EVAL_FIFO_DATA_WIDTH-1:0] neighbor_force_data_from_FIFO_2,
	input [NUM_PIPELINES-1:0] ref_force_valid,																// Meaning not empty
	input [NUM_PIPELINES-1:0] neighbor_force_valid_1,
	input [NUM_PIPELINES-1:0] neighbor_force_valid_2,
	input [CELL_ID_WIDTH-1:0] cellz,
	
	output [NUM_PIPELINES-1:0] ref_force_write_success,
	output [NUM_PIPELINES-1:0] neighbor_force_write_success_1,
	output [NUM_PIPELINES-1:0] neighbor_force_write_success_2, 
	output [TOTAL_CELL_NUM*FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values
);

reg [TOTAL_CELL_NUM*FORCE_EVAL_FIFO_DATA_WIDTH-1:0] reg_valid_force_values;
assign valid_force_values = reg_valid_force_values;

// Neighbor_1 mapping: 222, 223, 231, 232, 233, 311, 312 (LSB -> MSB)
// Neighbor_2 mapping: 313, 321, 322, 323, 331, 332, 333

wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_1_1_mid;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_1_2_mid;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_1_3_mid;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_1_4_mid;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_2_1_mid;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_2_2_mid;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_2_3_mid;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_2_4_mid;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_3_1_mid;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_3_2_mid;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_3_3_mid;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_3_4_mid;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_4_1_mid;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_4_2_mid;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_4_3_mid;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_4_4_mid;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_1_1_top;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_1_2_top;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_1_3_top;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_1_4_top;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_2_1_top;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_2_2_top;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_2_3_top;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_2_4_top;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_3_1_top;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_3_2_top;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_3_3_top;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_3_4_top;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_4_1_top;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_4_2_top;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_4_3_top;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_4_4_top;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_1_1_bottom;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_1_2_bottom;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_1_3_bottom;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_1_4_bottom;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_2_1_bottom;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_2_2_bottom;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_2_3_bottom;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_2_4_bottom;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_3_1_bottom;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_3_2_bottom;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_3_3_bottom;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_3_4_bottom;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_4_1_bottom;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_4_2_bottom;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_4_3_bottom;
wire [FORCE_WTADDR_ARBITER_SIZE-1:0] Arbitration_4_4_bottom;

assign ref_force_write_success[0] = Arbitration_1_1_mid[0];
assign ref_force_write_success[1] = Arbitration_1_2_mid[0];
assign ref_force_write_success[2] = Arbitration_1_3_mid[0];
assign ref_force_write_success[3] = Arbitration_1_4_mid[0];
assign ref_force_write_success[4] = Arbitration_2_1_mid[0];
assign ref_force_write_success[5] = Arbitration_2_2_mid[0];
assign ref_force_write_success[6] = Arbitration_2_3_mid[0];
assign ref_force_write_success[7] = Arbitration_2_4_mid[0];
assign ref_force_write_success[8] = Arbitration_3_1_mid[0];
assign ref_force_write_success[9] = Arbitration_3_2_mid[0];
assign ref_force_write_success[10] = Arbitration_3_3_mid[0];
assign ref_force_write_success[11] = Arbitration_3_4_mid[0];
assign ref_force_write_success[12] = Arbitration_4_1_mid[0];
assign ref_force_write_success[13] = Arbitration_4_2_mid[0];
assign ref_force_write_success[14] = Arbitration_4_3_mid[0];
assign ref_force_write_success[15] = Arbitration_4_4_mid[0];

assign neighbor_force_write_success_1[0] = Arbitration_1_1_mid[1] | Arbitration_1_1_top[1] | Arbitration_1_2_bottom[1] | Arbitration_1_2_mid[1] | Arbitration_1_2_top[1] | Arbitration_2_4_bottom[1] | Arbitration_2_4_mid[1];
assign neighbor_force_write_success_1[1] = Arbitration_1_2_mid[2] | Arbitration_1_2_top[2] | Arbitration_1_3_bottom[1] | Arbitration_1_3_mid[1] | Arbitration_1_3_top[1] | Arbitration_2_1_bottom[1] | Arbitration_2_1_mid[1];
assign neighbor_force_write_success_1[2] = Arbitration_1_3_mid[2] | Arbitration_1_3_top[2] | Arbitration_1_4_bottom[1] | Arbitration_1_4_mid[1] | Arbitration_1_4_top[1] | Arbitration_2_2_bottom[1] | Arbitration_2_2_mid[1];
assign neighbor_force_write_success_1[3] = Arbitration_1_4_mid[2] | Arbitration_1_4_top[2] | Arbitration_1_1_bottom[1] | Arbitration_1_1_mid[2] | Arbitration_1_1_top[2] | Arbitration_2_3_bottom[1] | Arbitration_2_3_mid[1];
assign neighbor_force_write_success_1[4] = Arbitration_2_1_mid[2] | Arbitration_2_1_top[1] | Arbitration_2_2_bottom[2] | Arbitration_2_2_mid[2] | Arbitration_2_2_top[1] | Arbitration_3_4_bottom[1] | Arbitration_3_4_mid[1];
assign neighbor_force_write_success_1[5] = Arbitration_2_2_mid[3] | Arbitration_2_2_top[2] | Arbitration_2_3_bottom[2] | Arbitration_2_3_mid[2] | Arbitration_2_3_top[1] | Arbitration_3_1_bottom[1] | Arbitration_3_1_mid[1];
assign neighbor_force_write_success_1[6] = Arbitration_2_3_mid[3] | Arbitration_2_3_top[2] | Arbitration_2_4_bottom[2] | Arbitration_2_4_mid[2] | Arbitration_2_4_top[1] | Arbitration_3_2_bottom[1] | Arbitration_3_2_mid[1];
assign neighbor_force_write_success_1[7] = Arbitration_2_4_mid[3] | Arbitration_2_4_top[2] | Arbitration_2_1_bottom[2] | Arbitration_2_1_mid[3] | Arbitration_2_1_top[2] | Arbitration_3_3_bottom[1] | Arbitration_3_3_mid[1];
assign neighbor_force_write_success_1[8] = Arbitration_3_1_mid[2] | Arbitration_3_1_top[1] | Arbitration_3_2_bottom[2] | Arbitration_3_2_mid[2] | Arbitration_3_2_top[1] | Arbitration_4_4_bottom[1] | Arbitration_4_4_mid[1];
assign neighbor_force_write_success_1[9] = Arbitration_3_2_mid[3] | Arbitration_3_2_top[2] | Arbitration_3_3_bottom[2] | Arbitration_3_3_mid[2] | Arbitration_3_3_top[1] | Arbitration_4_1_bottom[1] | Arbitration_4_1_mid[1];
assign neighbor_force_write_success_1[10] = Arbitration_3_3_mid[3] | Arbitration_3_3_top[2] | Arbitration_3_4_bottom[2] | Arbitration_3_4_mid[2] | Arbitration_3_4_top[1] | Arbitration_4_2_bottom[1] | Arbitration_4_2_mid[1];
assign neighbor_force_write_success_1[11] = Arbitration_3_4_mid[3] | Arbitration_3_4_top[2] | Arbitration_3_1_bottom[2] | Arbitration_3_1_mid[3] | Arbitration_3_1_top[2] | Arbitration_4_3_bottom[1] | Arbitration_4_3_mid[1];
assign neighbor_force_write_success_1[12] = Arbitration_4_1_mid[2] | Arbitration_4_1_top[1] | Arbitration_4_2_bottom[2] | Arbitration_4_2_mid[2] | Arbitration_4_2_top[1] | Arbitration_1_4_bottom[2] | Arbitration_1_4_mid[3];
assign neighbor_force_write_success_1[13] = Arbitration_4_2_mid[3] | Arbitration_4_2_top[2] | Arbitration_4_3_bottom[2] | Arbitration_4_3_mid[2] | Arbitration_4_3_top[1] | Arbitration_1_1_bottom[2] | Arbitration_1_1_mid[3];
assign neighbor_force_write_success_1[14] = Arbitration_4_3_mid[3] | Arbitration_4_3_top[2] | Arbitration_4_4_bottom[2] | Arbitration_4_4_mid[2] | Arbitration_4_4_top[1] | Arbitration_1_2_bottom[2] | Arbitration_1_2_mid[3];
assign neighbor_force_write_success_1[15] = Arbitration_4_4_mid[3] | Arbitration_4_4_top[2] | Arbitration_4_1_bottom[2] | Arbitration_4_1_mid[3] | Arbitration_4_1_top[2] | Arbitration_1_3_bottom[2] | Arbitration_1_3_mid[3];
assign neighbor_force_write_success_2[0] = Arbitration_2_4_top[3] | Arbitration_2_1_bottom[3] | Arbitration_2_1_mid[4] | Arbitration_2_1_top[3] | Arbitration_2_2_bottom[3] | Arbitration_2_2_mid[4] | Arbitration_2_2_top[3];
assign neighbor_force_write_success_2[1] = Arbitration_2_1_top[4] | Arbitration_2_2_bottom[4] | Arbitration_2_2_mid[5] | Arbitration_2_2_top[4] | Arbitration_2_3_bottom[3] | Arbitration_2_3_mid[4] | Arbitration_2_3_top[3];
assign neighbor_force_write_success_2[2] = Arbitration_2_2_top[5] | Arbitration_2_3_bottom[4] | Arbitration_2_3_mid[5] | Arbitration_2_3_top[4] | Arbitration_2_4_bottom[3] | Arbitration_2_4_mid[4] | Arbitration_2_4_top[4];
assign neighbor_force_write_success_2[3] = Arbitration_2_3_top[5] | Arbitration_2_4_bottom[4] | Arbitration_2_4_mid[5] | Arbitration_2_4_top[5] | Arbitration_2_1_bottom[4] | Arbitration_2_1_mid[5] | Arbitration_2_1_top[5];
assign neighbor_force_write_success_2[4] = Arbitration_3_4_top[3] | Arbitration_3_1_bottom[3] | Arbitration_3_1_mid[4] | Arbitration_3_1_top[3] | Arbitration_3_2_bottom[3] | Arbitration_3_2_mid[4] | Arbitration_3_2_top[3];
assign neighbor_force_write_success_2[5] = Arbitration_3_1_top[4] | Arbitration_3_2_bottom[4] | Arbitration_3_2_mid[5] | Arbitration_3_2_top[4] | Arbitration_3_3_bottom[3] | Arbitration_3_3_mid[4] | Arbitration_3_3_top[3];
assign neighbor_force_write_success_2[6] = Arbitration_3_2_top[5] | Arbitration_3_3_bottom[4] | Arbitration_3_3_mid[5] | Arbitration_3_3_top[4] | Arbitration_3_4_bottom[3] | Arbitration_3_4_mid[4] | Arbitration_3_4_top[4];
assign neighbor_force_write_success_2[7] = Arbitration_3_3_top[5] | Arbitration_3_4_bottom[4] | Arbitration_3_4_mid[5] | Arbitration_3_4_top[5] | Arbitration_3_1_bottom[4] | Arbitration_3_1_mid[5] | Arbitration_3_1_top[5];
assign neighbor_force_write_success_2[8] = Arbitration_4_4_top[3] | Arbitration_4_1_bottom[3] | Arbitration_4_1_mid[4] | Arbitration_4_1_top[3] | Arbitration_4_2_bottom[3] | Arbitration_4_2_mid[4] | Arbitration_4_2_top[3];
assign neighbor_force_write_success_2[9] = Arbitration_4_1_top[4] | Arbitration_4_2_bottom[4] | Arbitration_4_2_mid[5] | Arbitration_4_2_top[4] | Arbitration_4_3_bottom[3] | Arbitration_4_3_mid[4] | Arbitration_4_3_top[3];
assign neighbor_force_write_success_2[10] = Arbitration_4_2_top[5] | Arbitration_4_3_bottom[4] | Arbitration_4_3_mid[5] | Arbitration_4_3_top[4] | Arbitration_4_4_bottom[3] | Arbitration_4_4_mid[4] | Arbitration_4_4_top[4];
assign neighbor_force_write_success_2[11] = Arbitration_4_3_top[5] | Arbitration_4_4_bottom[4] | Arbitration_4_4_mid[5] | Arbitration_4_4_top[5] | Arbitration_4_1_bottom[4] | Arbitration_4_1_mid[5] | Arbitration_4_1_top[5];
assign neighbor_force_write_success_2[12] = Arbitration_1_4_top[3] | Arbitration_1_1_bottom[3] | Arbitration_1_1_mid[4] | Arbitration_1_1_top[3] | Arbitration_1_2_bottom[3] | Arbitration_1_2_mid[4] | Arbitration_1_2_top[3];
assign neighbor_force_write_success_2[13] = Arbitration_1_1_top[4] | Arbitration_1_2_bottom[4] | Arbitration_1_2_mid[5] | Arbitration_1_2_top[4] | Arbitration_1_3_bottom[3] | Arbitration_1_3_mid[4] | Arbitration_1_3_top[3];
assign neighbor_force_write_success_2[14] = Arbitration_1_2_top[5] | Arbitration_1_3_bottom[4] | Arbitration_1_3_mid[5] | Arbitration_1_3_top[4] | Arbitration_1_4_bottom[3] | Arbitration_1_4_mid[4] | Arbitration_1_4_top[4];
assign neighbor_force_write_success_2[15] = Arbitration_1_3_top[5] | Arbitration_1_4_bottom[4] | Arbitration_1_4_mid[5] | Arbitration_1_4_top[5] | Arbitration_1_1_bottom[4] | Arbitration_1_1_mid[5] | Arbitration_1_1_top[5];

reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_1_1_mid;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_1_2_mid;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_1_3_mid;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_1_4_mid;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_2_1_mid;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_2_2_mid;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_2_3_mid;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_2_4_mid;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_3_1_mid;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_3_2_mid;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_3_3_mid;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_3_4_mid;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_4_1_mid;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_4_2_mid;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_4_3_mid;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_4_4_mid;

reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_1_1_top;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_1_2_top;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_1_3_top;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_1_4_top;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_2_1_top;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_2_2_top;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_2_3_top;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_2_4_top;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_3_1_top;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_3_2_top;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_3_3_top;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_3_4_top;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_4_1_top;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_4_2_top;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_4_3_top;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_4_4_top;

reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_1_1_bottom;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_1_2_bottom;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_1_3_bottom;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_1_4_bottom;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_2_1_bottom;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_2_2_bottom;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_2_3_bottom;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_2_4_bottom;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_3_1_bottom;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_3_2_bottom;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_3_3_bottom;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_3_4_bottom;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_4_1_bottom;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_4_2_bottom;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_4_3_bottom;
reg [FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values_4_4_bottom;

reg force_valid_1_1_mid_1;
reg force_valid_1_1_mid_2;
reg force_valid_1_1_mid_3;
reg force_valid_1_1_mid_4;
reg force_valid_1_1_mid_5;
reg force_valid_1_1_top_1;
reg force_valid_1_1_top_2;
reg force_valid_1_1_top_3;
reg force_valid_1_1_top_4;
reg force_valid_1_1_top_5;
reg force_valid_1_1_bottom_1;
reg force_valid_1_1_bottom_2;
reg force_valid_1_1_bottom_3;
reg force_valid_1_1_bottom_4;
reg force_valid_1_1_bottom_5;
reg force_valid_1_2_mid_1;
reg force_valid_1_2_mid_2;
reg force_valid_1_2_mid_3;
reg force_valid_1_2_mid_4;
reg force_valid_1_2_mid_5;
reg force_valid_1_2_top_1;
reg force_valid_1_2_top_2;
reg force_valid_1_2_top_3;
reg force_valid_1_2_top_4;
reg force_valid_1_2_top_5;
reg force_valid_1_2_bottom_1;
reg force_valid_1_2_bottom_2;
reg force_valid_1_2_bottom_3;
reg force_valid_1_2_bottom_4;
reg force_valid_1_2_bottom_5;
reg force_valid_1_3_mid_1;
reg force_valid_1_3_mid_2;
reg force_valid_1_3_mid_3;
reg force_valid_1_3_mid_4;
reg force_valid_1_3_mid_5;
reg force_valid_1_3_top_1;
reg force_valid_1_3_top_2;
reg force_valid_1_3_top_3;
reg force_valid_1_3_top_4;
reg force_valid_1_3_top_5;
reg force_valid_1_3_bottom_1;
reg force_valid_1_3_bottom_2;
reg force_valid_1_3_bottom_3;
reg force_valid_1_3_bottom_4;
reg force_valid_1_3_bottom_5;
reg force_valid_1_4_mid_1;
reg force_valid_1_4_mid_2;
reg force_valid_1_4_mid_3;
reg force_valid_1_4_mid_4;
reg force_valid_1_4_mid_5;
reg force_valid_1_4_top_1;
reg force_valid_1_4_top_2;
reg force_valid_1_4_top_3;
reg force_valid_1_4_top_4;
reg force_valid_1_4_top_5;
reg force_valid_1_4_bottom_1;
reg force_valid_1_4_bottom_2;
reg force_valid_1_4_bottom_3;
reg force_valid_1_4_bottom_4;
reg force_valid_1_4_bottom_5;
reg force_valid_2_1_mid_1;
reg force_valid_2_1_mid_2;
reg force_valid_2_1_mid_3;
reg force_valid_2_1_mid_4;
reg force_valid_2_1_mid_5;
reg force_valid_2_1_top_1;
reg force_valid_2_1_top_2;
reg force_valid_2_1_top_3;
reg force_valid_2_1_top_4;
reg force_valid_2_1_top_5;
reg force_valid_2_1_bottom_1;
reg force_valid_2_1_bottom_2;
reg force_valid_2_1_bottom_3;
reg force_valid_2_1_bottom_4;
reg force_valid_2_1_bottom_5;
reg force_valid_2_2_mid_1;
reg force_valid_2_2_mid_2;
reg force_valid_2_2_mid_3;
reg force_valid_2_2_mid_4;
reg force_valid_2_2_mid_5;
reg force_valid_2_2_top_1;
reg force_valid_2_2_top_2;
reg force_valid_2_2_top_3;
reg force_valid_2_2_top_4;
reg force_valid_2_2_top_5;
reg force_valid_2_2_bottom_1;
reg force_valid_2_2_bottom_2;
reg force_valid_2_2_bottom_3;
reg force_valid_2_2_bottom_4;
reg force_valid_2_2_bottom_5;
reg force_valid_2_3_mid_1;
reg force_valid_2_3_mid_2;
reg force_valid_2_3_mid_3;
reg force_valid_2_3_mid_4;
reg force_valid_2_3_mid_5;
reg force_valid_2_3_top_1;
reg force_valid_2_3_top_2;
reg force_valid_2_3_top_3;
reg force_valid_2_3_top_4;
reg force_valid_2_3_top_5;
reg force_valid_2_3_bottom_1;
reg force_valid_2_3_bottom_2;
reg force_valid_2_3_bottom_3;
reg force_valid_2_3_bottom_4;
reg force_valid_2_3_bottom_5;
reg force_valid_2_4_mid_1;
reg force_valid_2_4_mid_2;
reg force_valid_2_4_mid_3;
reg force_valid_2_4_mid_4;
reg force_valid_2_4_mid_5;
reg force_valid_2_4_top_1;
reg force_valid_2_4_top_2;
reg force_valid_2_4_top_3;
reg force_valid_2_4_top_4;
reg force_valid_2_4_top_5;
reg force_valid_2_4_bottom_1;
reg force_valid_2_4_bottom_2;
reg force_valid_2_4_bottom_3;
reg force_valid_2_4_bottom_4;
reg force_valid_2_4_bottom_5;
reg force_valid_3_1_mid_1;
reg force_valid_3_1_mid_2;
reg force_valid_3_1_mid_3;
reg force_valid_3_1_mid_4;
reg force_valid_3_1_mid_5;
reg force_valid_3_1_top_1;
reg force_valid_3_1_top_2;
reg force_valid_3_1_top_3;
reg force_valid_3_1_top_4;
reg force_valid_3_1_top_5;
reg force_valid_3_1_bottom_1;
reg force_valid_3_1_bottom_2;
reg force_valid_3_1_bottom_3;
reg force_valid_3_1_bottom_4;
reg force_valid_3_1_bottom_5;
reg force_valid_3_2_mid_1;
reg force_valid_3_2_mid_2;
reg force_valid_3_2_mid_3;
reg force_valid_3_2_mid_4;
reg force_valid_3_2_mid_5;
reg force_valid_3_2_top_1;
reg force_valid_3_2_top_2;
reg force_valid_3_2_top_3;
reg force_valid_3_2_top_4;
reg force_valid_3_2_top_5;
reg force_valid_3_2_bottom_1;
reg force_valid_3_2_bottom_2;
reg force_valid_3_2_bottom_3;
reg force_valid_3_2_bottom_4;
reg force_valid_3_2_bottom_5;
reg force_valid_3_3_mid_1;
reg force_valid_3_3_mid_2;
reg force_valid_3_3_mid_3;
reg force_valid_3_3_mid_4;
reg force_valid_3_3_mid_5;
reg force_valid_3_3_top_1;
reg force_valid_3_3_top_2;
reg force_valid_3_3_top_3;
reg force_valid_3_3_top_4;
reg force_valid_3_3_top_5;
reg force_valid_3_3_bottom_1;
reg force_valid_3_3_bottom_2;
reg force_valid_3_3_bottom_3;
reg force_valid_3_3_bottom_4;
reg force_valid_3_3_bottom_5;
reg force_valid_3_4_mid_1;
reg force_valid_3_4_mid_2;
reg force_valid_3_4_mid_3;
reg force_valid_3_4_mid_4;
reg force_valid_3_4_mid_5;
reg force_valid_3_4_top_1;
reg force_valid_3_4_top_2;
reg force_valid_3_4_top_3;
reg force_valid_3_4_top_4;
reg force_valid_3_4_top_5;
reg force_valid_3_4_bottom_1;
reg force_valid_3_4_bottom_2;
reg force_valid_3_4_bottom_3;
reg force_valid_3_4_bottom_4;
reg force_valid_3_4_bottom_5;
reg force_valid_4_1_mid_1;
reg force_valid_4_1_mid_2;
reg force_valid_4_1_mid_3;
reg force_valid_4_1_mid_4;
reg force_valid_4_1_mid_5;
reg force_valid_4_1_top_1;
reg force_valid_4_1_top_2;
reg force_valid_4_1_top_3;
reg force_valid_4_1_top_4;
reg force_valid_4_1_top_5;
reg force_valid_4_1_bottom_1;
reg force_valid_4_1_bottom_2;
reg force_valid_4_1_bottom_3;
reg force_valid_4_1_bottom_4;
reg force_valid_4_1_bottom_5;
reg force_valid_4_2_mid_1;
reg force_valid_4_2_mid_2;
reg force_valid_4_2_mid_3;
reg force_valid_4_2_mid_4;
reg force_valid_4_2_mid_5;
reg force_valid_4_2_top_1;
reg force_valid_4_2_top_2;
reg force_valid_4_2_top_3;
reg force_valid_4_2_top_4;
reg force_valid_4_2_top_5;
reg force_valid_4_2_bottom_1;
reg force_valid_4_2_bottom_2;
reg force_valid_4_2_bottom_3;
reg force_valid_4_2_bottom_4;
reg force_valid_4_2_bottom_5;
reg force_valid_4_3_mid_1;
reg force_valid_4_3_mid_2;
reg force_valid_4_3_mid_3;
reg force_valid_4_3_mid_4;
reg force_valid_4_3_mid_5;
reg force_valid_4_3_top_1;
reg force_valid_4_3_top_2;
reg force_valid_4_3_top_3;
reg force_valid_4_3_top_4;
reg force_valid_4_3_top_5;
reg force_valid_4_3_bottom_1;
reg force_valid_4_3_bottom_2;
reg force_valid_4_3_bottom_3;
reg force_valid_4_3_bottom_4;
reg force_valid_4_3_bottom_5;
reg force_valid_4_4_mid_1;
reg force_valid_4_4_mid_2;
reg force_valid_4_4_mid_3;
reg force_valid_4_4_mid_4;
reg force_valid_4_4_mid_5;
reg force_valid_4_4_top_1;
reg force_valid_4_4_top_2;
reg force_valid_4_4_top_3;
reg force_valid_4_4_top_4;
reg force_valid_4_4_top_5;
reg force_valid_4_4_bottom_1;
reg force_valid_4_4_bottom_2;
reg force_valid_4_4_bottom_3;
reg force_valid_4_4_bottom_4;
reg force_valid_4_4_bottom_5;
always@(*)
	begin
	case(cellz)
		1:
			begin
			reg_valid_force_values[3*FORCE_EVAL_FIFO_DATA_WIDTH-1:2*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[7*FORCE_EVAL_FIFO_DATA_WIDTH-1:6*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[11*FORCE_EVAL_FIFO_DATA_WIDTH-1:10*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[15*FORCE_EVAL_FIFO_DATA_WIDTH-1:14*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[19*FORCE_EVAL_FIFO_DATA_WIDTH-1:18*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[23*FORCE_EVAL_FIFO_DATA_WIDTH-1:22*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[27*FORCE_EVAL_FIFO_DATA_WIDTH-1:26*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[31*FORCE_EVAL_FIFO_DATA_WIDTH-1:30*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[35*FORCE_EVAL_FIFO_DATA_WIDTH-1:34*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[39*FORCE_EVAL_FIFO_DATA_WIDTH-1:38*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[43*FORCE_EVAL_FIFO_DATA_WIDTH-1:42*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[47*FORCE_EVAL_FIFO_DATA_WIDTH-1:46*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[51*FORCE_EVAL_FIFO_DATA_WIDTH-1:50*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[55*FORCE_EVAL_FIFO_DATA_WIDTH-1:54*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[59*FORCE_EVAL_FIFO_DATA_WIDTH-1:58*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[63*FORCE_EVAL_FIFO_DATA_WIDTH-1:62*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[1*FORCE_EVAL_FIFO_DATA_WIDTH-1:0*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_1_mid;
			reg_valid_force_values[2*FORCE_EVAL_FIFO_DATA_WIDTH-1:1*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_1_top;
			reg_valid_force_values[4*FORCE_EVAL_FIFO_DATA_WIDTH-1:3*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_1_bottom;
			reg_valid_force_values[5*FORCE_EVAL_FIFO_DATA_WIDTH-1:4*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_2_mid;
			reg_valid_force_values[6*FORCE_EVAL_FIFO_DATA_WIDTH-1:5*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_2_top;
			reg_valid_force_values[8*FORCE_EVAL_FIFO_DATA_WIDTH-1:7*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_2_bottom;
			reg_valid_force_values[9*FORCE_EVAL_FIFO_DATA_WIDTH-1:8*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_3_mid;
			reg_valid_force_values[10*FORCE_EVAL_FIFO_DATA_WIDTH-1:9*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_3_top;
			reg_valid_force_values[12*FORCE_EVAL_FIFO_DATA_WIDTH-1:11*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_3_bottom;
			reg_valid_force_values[13*FORCE_EVAL_FIFO_DATA_WIDTH-1:12*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_4_mid;
			reg_valid_force_values[14*FORCE_EVAL_FIFO_DATA_WIDTH-1:13*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_4_top;
			reg_valid_force_values[16*FORCE_EVAL_FIFO_DATA_WIDTH-1:15*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_4_bottom;
			reg_valid_force_values[17*FORCE_EVAL_FIFO_DATA_WIDTH-1:16*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_1_mid;
			reg_valid_force_values[18*FORCE_EVAL_FIFO_DATA_WIDTH-1:17*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_1_top;
			reg_valid_force_values[20*FORCE_EVAL_FIFO_DATA_WIDTH-1:19*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_1_bottom;
			reg_valid_force_values[21*FORCE_EVAL_FIFO_DATA_WIDTH-1:20*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_2_mid;
			reg_valid_force_values[22*FORCE_EVAL_FIFO_DATA_WIDTH-1:21*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_2_top;
			reg_valid_force_values[24*FORCE_EVAL_FIFO_DATA_WIDTH-1:23*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_2_bottom;
			reg_valid_force_values[25*FORCE_EVAL_FIFO_DATA_WIDTH-1:24*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_3_mid;
			reg_valid_force_values[26*FORCE_EVAL_FIFO_DATA_WIDTH-1:25*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_3_top;
			reg_valid_force_values[28*FORCE_EVAL_FIFO_DATA_WIDTH-1:27*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_3_bottom;
			reg_valid_force_values[29*FORCE_EVAL_FIFO_DATA_WIDTH-1:28*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_4_mid;
			reg_valid_force_values[30*FORCE_EVAL_FIFO_DATA_WIDTH-1:29*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_4_top;
			reg_valid_force_values[32*FORCE_EVAL_FIFO_DATA_WIDTH-1:31*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_4_bottom;
			reg_valid_force_values[33*FORCE_EVAL_FIFO_DATA_WIDTH-1:32*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_1_mid;
			reg_valid_force_values[34*FORCE_EVAL_FIFO_DATA_WIDTH-1:33*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_1_top;
			reg_valid_force_values[36*FORCE_EVAL_FIFO_DATA_WIDTH-1:35*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_1_bottom;
			reg_valid_force_values[37*FORCE_EVAL_FIFO_DATA_WIDTH-1:36*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_2_mid;
			reg_valid_force_values[38*FORCE_EVAL_FIFO_DATA_WIDTH-1:37*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_2_top;
			reg_valid_force_values[40*FORCE_EVAL_FIFO_DATA_WIDTH-1:39*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_2_bottom;
			reg_valid_force_values[41*FORCE_EVAL_FIFO_DATA_WIDTH-1:40*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_3_mid;
			reg_valid_force_values[42*FORCE_EVAL_FIFO_DATA_WIDTH-1:41*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_3_top;
			reg_valid_force_values[44*FORCE_EVAL_FIFO_DATA_WIDTH-1:43*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_3_bottom;
			reg_valid_force_values[45*FORCE_EVAL_FIFO_DATA_WIDTH-1:44*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_4_mid;
			reg_valid_force_values[46*FORCE_EVAL_FIFO_DATA_WIDTH-1:45*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_4_top;
			reg_valid_force_values[48*FORCE_EVAL_FIFO_DATA_WIDTH-1:47*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_4_bottom;
			reg_valid_force_values[49*FORCE_EVAL_FIFO_DATA_WIDTH-1:48*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_1_mid;
			reg_valid_force_values[50*FORCE_EVAL_FIFO_DATA_WIDTH-1:49*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_1_top;
			reg_valid_force_values[52*FORCE_EVAL_FIFO_DATA_WIDTH-1:51*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_1_bottom;
			reg_valid_force_values[53*FORCE_EVAL_FIFO_DATA_WIDTH-1:52*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_2_mid;
			reg_valid_force_values[54*FORCE_EVAL_FIFO_DATA_WIDTH-1:53*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_2_top;
			reg_valid_force_values[56*FORCE_EVAL_FIFO_DATA_WIDTH-1:55*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_2_bottom;
			reg_valid_force_values[57*FORCE_EVAL_FIFO_DATA_WIDTH-1:56*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_3_mid;
			reg_valid_force_values[58*FORCE_EVAL_FIFO_DATA_WIDTH-1:57*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_3_top;
			reg_valid_force_values[60*FORCE_EVAL_FIFO_DATA_WIDTH-1:59*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_3_bottom;
			reg_valid_force_values[61*FORCE_EVAL_FIFO_DATA_WIDTH-1:60*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_4_mid;
			reg_valid_force_values[62*FORCE_EVAL_FIFO_DATA_WIDTH-1:61*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_4_top;
			reg_valid_force_values[64*FORCE_EVAL_FIFO_DATA_WIDTH-1:63*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_4_bottom;
			end
		2:
			begin
			reg_valid_force_values[4*FORCE_EVAL_FIFO_DATA_WIDTH-1:3*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[8*FORCE_EVAL_FIFO_DATA_WIDTH-1:7*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[12*FORCE_EVAL_FIFO_DATA_WIDTH-1:11*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[16*FORCE_EVAL_FIFO_DATA_WIDTH-1:15*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[20*FORCE_EVAL_FIFO_DATA_WIDTH-1:19*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[24*FORCE_EVAL_FIFO_DATA_WIDTH-1:23*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[28*FORCE_EVAL_FIFO_DATA_WIDTH-1:27*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[32*FORCE_EVAL_FIFO_DATA_WIDTH-1:31*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[36*FORCE_EVAL_FIFO_DATA_WIDTH-1:35*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[40*FORCE_EVAL_FIFO_DATA_WIDTH-1:39*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[44*FORCE_EVAL_FIFO_DATA_WIDTH-1:43*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[48*FORCE_EVAL_FIFO_DATA_WIDTH-1:47*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[52*FORCE_EVAL_FIFO_DATA_WIDTH-1:51*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[56*FORCE_EVAL_FIFO_DATA_WIDTH-1:55*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[60*FORCE_EVAL_FIFO_DATA_WIDTH-1:59*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[64*FORCE_EVAL_FIFO_DATA_WIDTH-1:63*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[2*FORCE_EVAL_FIFO_DATA_WIDTH-1:1*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_1_mid;
			reg_valid_force_values[3*FORCE_EVAL_FIFO_DATA_WIDTH-1:2*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_1_top;
			reg_valid_force_values[1*FORCE_EVAL_FIFO_DATA_WIDTH-1:0*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_1_bottom;
			reg_valid_force_values[6*FORCE_EVAL_FIFO_DATA_WIDTH-1:5*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_2_mid;
			reg_valid_force_values[7*FORCE_EVAL_FIFO_DATA_WIDTH-1:6*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_2_top;
			reg_valid_force_values[5*FORCE_EVAL_FIFO_DATA_WIDTH-1:4*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_2_bottom;
			reg_valid_force_values[10*FORCE_EVAL_FIFO_DATA_WIDTH-1:9*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_3_mid;
			reg_valid_force_values[11*FORCE_EVAL_FIFO_DATA_WIDTH-1:10*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_3_top;
			reg_valid_force_values[9*FORCE_EVAL_FIFO_DATA_WIDTH-1:8*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_3_bottom;
			reg_valid_force_values[14*FORCE_EVAL_FIFO_DATA_WIDTH-1:13*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_4_mid;
			reg_valid_force_values[15*FORCE_EVAL_FIFO_DATA_WIDTH-1:14*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_4_top;
			reg_valid_force_values[13*FORCE_EVAL_FIFO_DATA_WIDTH-1:12*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_4_bottom;
			reg_valid_force_values[18*FORCE_EVAL_FIFO_DATA_WIDTH-1:17*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_1_mid;
			reg_valid_force_values[19*FORCE_EVAL_FIFO_DATA_WIDTH-1:18*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_1_top;
			reg_valid_force_values[17*FORCE_EVAL_FIFO_DATA_WIDTH-1:16*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_1_bottom;
			reg_valid_force_values[22*FORCE_EVAL_FIFO_DATA_WIDTH-1:21*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_2_mid;
			reg_valid_force_values[23*FORCE_EVAL_FIFO_DATA_WIDTH-1:22*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_2_top;
			reg_valid_force_values[21*FORCE_EVAL_FIFO_DATA_WIDTH-1:20*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_2_bottom;
			reg_valid_force_values[26*FORCE_EVAL_FIFO_DATA_WIDTH-1:25*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_3_mid;
			reg_valid_force_values[27*FORCE_EVAL_FIFO_DATA_WIDTH-1:26*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_3_top;
			reg_valid_force_values[25*FORCE_EVAL_FIFO_DATA_WIDTH-1:24*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_3_bottom;
			reg_valid_force_values[30*FORCE_EVAL_FIFO_DATA_WIDTH-1:29*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_4_mid;
			reg_valid_force_values[31*FORCE_EVAL_FIFO_DATA_WIDTH-1:30*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_4_top;
			reg_valid_force_values[29*FORCE_EVAL_FIFO_DATA_WIDTH-1:28*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_4_bottom;
			reg_valid_force_values[34*FORCE_EVAL_FIFO_DATA_WIDTH-1:33*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_1_mid;
			reg_valid_force_values[35*FORCE_EVAL_FIFO_DATA_WIDTH-1:34*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_1_top;
			reg_valid_force_values[33*FORCE_EVAL_FIFO_DATA_WIDTH-1:32*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_1_bottom;
			reg_valid_force_values[38*FORCE_EVAL_FIFO_DATA_WIDTH-1:37*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_2_mid;
			reg_valid_force_values[39*FORCE_EVAL_FIFO_DATA_WIDTH-1:38*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_2_top;
			reg_valid_force_values[37*FORCE_EVAL_FIFO_DATA_WIDTH-1:36*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_2_bottom;
			reg_valid_force_values[42*FORCE_EVAL_FIFO_DATA_WIDTH-1:41*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_3_mid;
			reg_valid_force_values[43*FORCE_EVAL_FIFO_DATA_WIDTH-1:42*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_3_top;
			reg_valid_force_values[41*FORCE_EVAL_FIFO_DATA_WIDTH-1:40*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_3_bottom;
			reg_valid_force_values[46*FORCE_EVAL_FIFO_DATA_WIDTH-1:45*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_4_mid;
			reg_valid_force_values[47*FORCE_EVAL_FIFO_DATA_WIDTH-1:46*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_4_top;
			reg_valid_force_values[45*FORCE_EVAL_FIFO_DATA_WIDTH-1:44*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_4_bottom;
			reg_valid_force_values[50*FORCE_EVAL_FIFO_DATA_WIDTH-1:49*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_1_mid;
			reg_valid_force_values[51*FORCE_EVAL_FIFO_DATA_WIDTH-1:50*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_1_top;
			reg_valid_force_values[49*FORCE_EVAL_FIFO_DATA_WIDTH-1:48*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_1_bottom;
			reg_valid_force_values[54*FORCE_EVAL_FIFO_DATA_WIDTH-1:53*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_2_mid;
			reg_valid_force_values[55*FORCE_EVAL_FIFO_DATA_WIDTH-1:54*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_2_top;
			reg_valid_force_values[53*FORCE_EVAL_FIFO_DATA_WIDTH-1:52*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_2_bottom;
			reg_valid_force_values[58*FORCE_EVAL_FIFO_DATA_WIDTH-1:57*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_3_mid;
			reg_valid_force_values[59*FORCE_EVAL_FIFO_DATA_WIDTH-1:58*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_3_top;
			reg_valid_force_values[57*FORCE_EVAL_FIFO_DATA_WIDTH-1:56*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_3_bottom;
			reg_valid_force_values[62*FORCE_EVAL_FIFO_DATA_WIDTH-1:61*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_4_mid;
			reg_valid_force_values[63*FORCE_EVAL_FIFO_DATA_WIDTH-1:62*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_4_top;
			reg_valid_force_values[61*FORCE_EVAL_FIFO_DATA_WIDTH-1:60*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_4_bottom;
			end
		3:
			begin
			reg_valid_force_values[1*FORCE_EVAL_FIFO_DATA_WIDTH-1:0*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[5*FORCE_EVAL_FIFO_DATA_WIDTH-1:4*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[9*FORCE_EVAL_FIFO_DATA_WIDTH-1:8*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[13*FORCE_EVAL_FIFO_DATA_WIDTH-1:12*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[17*FORCE_EVAL_FIFO_DATA_WIDTH-1:16*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[21*FORCE_EVAL_FIFO_DATA_WIDTH-1:20*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[25*FORCE_EVAL_FIFO_DATA_WIDTH-1:24*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[29*FORCE_EVAL_FIFO_DATA_WIDTH-1:28*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[33*FORCE_EVAL_FIFO_DATA_WIDTH-1:32*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[37*FORCE_EVAL_FIFO_DATA_WIDTH-1:36*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[41*FORCE_EVAL_FIFO_DATA_WIDTH-1:40*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[45*FORCE_EVAL_FIFO_DATA_WIDTH-1:44*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[49*FORCE_EVAL_FIFO_DATA_WIDTH-1:48*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[53*FORCE_EVAL_FIFO_DATA_WIDTH-1:52*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[57*FORCE_EVAL_FIFO_DATA_WIDTH-1:56*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[61*FORCE_EVAL_FIFO_DATA_WIDTH-1:60*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[3*FORCE_EVAL_FIFO_DATA_WIDTH-1:2*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_1_mid;
			reg_valid_force_values[4*FORCE_EVAL_FIFO_DATA_WIDTH-1:3*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_1_top;
			reg_valid_force_values[2*FORCE_EVAL_FIFO_DATA_WIDTH-1:1*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_1_bottom;
			reg_valid_force_values[7*FORCE_EVAL_FIFO_DATA_WIDTH-1:6*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_2_mid;
			reg_valid_force_values[8*FORCE_EVAL_FIFO_DATA_WIDTH-1:7*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_2_top;
			reg_valid_force_values[6*FORCE_EVAL_FIFO_DATA_WIDTH-1:5*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_2_bottom;
			reg_valid_force_values[11*FORCE_EVAL_FIFO_DATA_WIDTH-1:10*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_3_mid;
			reg_valid_force_values[12*FORCE_EVAL_FIFO_DATA_WIDTH-1:11*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_3_top;
			reg_valid_force_values[10*FORCE_EVAL_FIFO_DATA_WIDTH-1:9*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_3_bottom;
			reg_valid_force_values[15*FORCE_EVAL_FIFO_DATA_WIDTH-1:14*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_4_mid;
			reg_valid_force_values[16*FORCE_EVAL_FIFO_DATA_WIDTH-1:15*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_4_top;
			reg_valid_force_values[14*FORCE_EVAL_FIFO_DATA_WIDTH-1:13*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_4_bottom;
			reg_valid_force_values[19*FORCE_EVAL_FIFO_DATA_WIDTH-1:18*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_1_mid;
			reg_valid_force_values[20*FORCE_EVAL_FIFO_DATA_WIDTH-1:19*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_1_top;
			reg_valid_force_values[18*FORCE_EVAL_FIFO_DATA_WIDTH-1:17*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_1_bottom;
			reg_valid_force_values[23*FORCE_EVAL_FIFO_DATA_WIDTH-1:22*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_2_mid;
			reg_valid_force_values[24*FORCE_EVAL_FIFO_DATA_WIDTH-1:23*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_2_top;
			reg_valid_force_values[22*FORCE_EVAL_FIFO_DATA_WIDTH-1:21*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_2_bottom;
			reg_valid_force_values[27*FORCE_EVAL_FIFO_DATA_WIDTH-1:26*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_3_mid;
			reg_valid_force_values[28*FORCE_EVAL_FIFO_DATA_WIDTH-1:27*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_3_top;
			reg_valid_force_values[26*FORCE_EVAL_FIFO_DATA_WIDTH-1:25*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_3_bottom;
			reg_valid_force_values[31*FORCE_EVAL_FIFO_DATA_WIDTH-1:30*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_4_mid;
			reg_valid_force_values[32*FORCE_EVAL_FIFO_DATA_WIDTH-1:31*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_4_top;
			reg_valid_force_values[30*FORCE_EVAL_FIFO_DATA_WIDTH-1:29*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_4_bottom;
			reg_valid_force_values[35*FORCE_EVAL_FIFO_DATA_WIDTH-1:34*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_1_mid;
			reg_valid_force_values[36*FORCE_EVAL_FIFO_DATA_WIDTH-1:35*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_1_top;
			reg_valid_force_values[34*FORCE_EVAL_FIFO_DATA_WIDTH-1:33*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_1_bottom;
			reg_valid_force_values[39*FORCE_EVAL_FIFO_DATA_WIDTH-1:38*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_2_mid;
			reg_valid_force_values[40*FORCE_EVAL_FIFO_DATA_WIDTH-1:39*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_2_top;
			reg_valid_force_values[38*FORCE_EVAL_FIFO_DATA_WIDTH-1:37*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_2_bottom;
			reg_valid_force_values[43*FORCE_EVAL_FIFO_DATA_WIDTH-1:42*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_3_mid;
			reg_valid_force_values[44*FORCE_EVAL_FIFO_DATA_WIDTH-1:43*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_3_top;
			reg_valid_force_values[42*FORCE_EVAL_FIFO_DATA_WIDTH-1:41*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_3_bottom;
			reg_valid_force_values[47*FORCE_EVAL_FIFO_DATA_WIDTH-1:46*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_4_mid;
			reg_valid_force_values[48*FORCE_EVAL_FIFO_DATA_WIDTH-1:47*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_4_top;
			reg_valid_force_values[46*FORCE_EVAL_FIFO_DATA_WIDTH-1:45*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_4_bottom;
			reg_valid_force_values[51*FORCE_EVAL_FIFO_DATA_WIDTH-1:50*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_1_mid;
			reg_valid_force_values[52*FORCE_EVAL_FIFO_DATA_WIDTH-1:51*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_1_top;
			reg_valid_force_values[50*FORCE_EVAL_FIFO_DATA_WIDTH-1:49*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_1_bottom;
			reg_valid_force_values[55*FORCE_EVAL_FIFO_DATA_WIDTH-1:54*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_2_mid;
			reg_valid_force_values[56*FORCE_EVAL_FIFO_DATA_WIDTH-1:55*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_2_top;
			reg_valid_force_values[54*FORCE_EVAL_FIFO_DATA_WIDTH-1:53*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_2_bottom;
			reg_valid_force_values[59*FORCE_EVAL_FIFO_DATA_WIDTH-1:58*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_3_mid;
			reg_valid_force_values[60*FORCE_EVAL_FIFO_DATA_WIDTH-1:59*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_3_top;
			reg_valid_force_values[58*FORCE_EVAL_FIFO_DATA_WIDTH-1:57*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_3_bottom;
			reg_valid_force_values[63*FORCE_EVAL_FIFO_DATA_WIDTH-1:62*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_4_mid;
			reg_valid_force_values[64*FORCE_EVAL_FIFO_DATA_WIDTH-1:63*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_4_top;
			reg_valid_force_values[62*FORCE_EVAL_FIFO_DATA_WIDTH-1:61*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_4_bottom;
			end
		4:
			begin
			reg_valid_force_values[2*FORCE_EVAL_FIFO_DATA_WIDTH-1:1*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[6*FORCE_EVAL_FIFO_DATA_WIDTH-1:5*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[10*FORCE_EVAL_FIFO_DATA_WIDTH-1:9*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[14*FORCE_EVAL_FIFO_DATA_WIDTH-1:13*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[18*FORCE_EVAL_FIFO_DATA_WIDTH-1:17*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[22*FORCE_EVAL_FIFO_DATA_WIDTH-1:21*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[26*FORCE_EVAL_FIFO_DATA_WIDTH-1:25*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[30*FORCE_EVAL_FIFO_DATA_WIDTH-1:29*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[34*FORCE_EVAL_FIFO_DATA_WIDTH-1:33*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[38*FORCE_EVAL_FIFO_DATA_WIDTH-1:37*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[42*FORCE_EVAL_FIFO_DATA_WIDTH-1:41*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[46*FORCE_EVAL_FIFO_DATA_WIDTH-1:45*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[50*FORCE_EVAL_FIFO_DATA_WIDTH-1:49*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[54*FORCE_EVAL_FIFO_DATA_WIDTH-1:53*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[58*FORCE_EVAL_FIFO_DATA_WIDTH-1:57*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[62*FORCE_EVAL_FIFO_DATA_WIDTH-1:61*FORCE_EVAL_FIFO_DATA_WIDTH] = 0;
			reg_valid_force_values[4*FORCE_EVAL_FIFO_DATA_WIDTH-1:3*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_1_mid;
			reg_valid_force_values[1*FORCE_EVAL_FIFO_DATA_WIDTH-1:0*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_1_top;
			reg_valid_force_values[3*FORCE_EVAL_FIFO_DATA_WIDTH-1:2*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_1_bottom;
			reg_valid_force_values[8*FORCE_EVAL_FIFO_DATA_WIDTH-1:7*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_2_mid;
			reg_valid_force_values[5*FORCE_EVAL_FIFO_DATA_WIDTH-1:4*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_2_top;
			reg_valid_force_values[7*FORCE_EVAL_FIFO_DATA_WIDTH-1:6*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_2_bottom;
			reg_valid_force_values[12*FORCE_EVAL_FIFO_DATA_WIDTH-1:11*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_3_mid;
			reg_valid_force_values[9*FORCE_EVAL_FIFO_DATA_WIDTH-1:8*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_3_top;
			reg_valid_force_values[11*FORCE_EVAL_FIFO_DATA_WIDTH-1:10*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_3_bottom;
			reg_valid_force_values[16*FORCE_EVAL_FIFO_DATA_WIDTH-1:15*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_4_mid;
			reg_valid_force_values[13*FORCE_EVAL_FIFO_DATA_WIDTH-1:12*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_4_top;
			reg_valid_force_values[15*FORCE_EVAL_FIFO_DATA_WIDTH-1:14*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_1_4_bottom;
			reg_valid_force_values[20*FORCE_EVAL_FIFO_DATA_WIDTH-1:19*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_1_mid;
			reg_valid_force_values[17*FORCE_EVAL_FIFO_DATA_WIDTH-1:16*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_1_top;
			reg_valid_force_values[19*FORCE_EVAL_FIFO_DATA_WIDTH-1:18*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_1_bottom;
			reg_valid_force_values[24*FORCE_EVAL_FIFO_DATA_WIDTH-1:23*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_2_mid;
			reg_valid_force_values[21*FORCE_EVAL_FIFO_DATA_WIDTH-1:20*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_2_top;
			reg_valid_force_values[23*FORCE_EVAL_FIFO_DATA_WIDTH-1:22*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_2_bottom;
			reg_valid_force_values[28*FORCE_EVAL_FIFO_DATA_WIDTH-1:27*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_3_mid;
			reg_valid_force_values[25*FORCE_EVAL_FIFO_DATA_WIDTH-1:24*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_3_top;
			reg_valid_force_values[27*FORCE_EVAL_FIFO_DATA_WIDTH-1:26*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_3_bottom;
			reg_valid_force_values[32*FORCE_EVAL_FIFO_DATA_WIDTH-1:31*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_4_mid;
			reg_valid_force_values[29*FORCE_EVAL_FIFO_DATA_WIDTH-1:28*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_4_top;
			reg_valid_force_values[31*FORCE_EVAL_FIFO_DATA_WIDTH-1:30*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_2_4_bottom;
			reg_valid_force_values[36*FORCE_EVAL_FIFO_DATA_WIDTH-1:35*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_1_mid;
			reg_valid_force_values[33*FORCE_EVAL_FIFO_DATA_WIDTH-1:32*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_1_top;
			reg_valid_force_values[35*FORCE_EVAL_FIFO_DATA_WIDTH-1:34*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_1_bottom;
			reg_valid_force_values[40*FORCE_EVAL_FIFO_DATA_WIDTH-1:39*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_2_mid;
			reg_valid_force_values[37*FORCE_EVAL_FIFO_DATA_WIDTH-1:36*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_2_top;
			reg_valid_force_values[39*FORCE_EVAL_FIFO_DATA_WIDTH-1:38*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_2_bottom;
			reg_valid_force_values[44*FORCE_EVAL_FIFO_DATA_WIDTH-1:43*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_3_mid;
			reg_valid_force_values[41*FORCE_EVAL_FIFO_DATA_WIDTH-1:40*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_3_top;
			reg_valid_force_values[43*FORCE_EVAL_FIFO_DATA_WIDTH-1:42*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_3_bottom;
			reg_valid_force_values[48*FORCE_EVAL_FIFO_DATA_WIDTH-1:47*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_4_mid;
			reg_valid_force_values[45*FORCE_EVAL_FIFO_DATA_WIDTH-1:44*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_4_top;
			reg_valid_force_values[47*FORCE_EVAL_FIFO_DATA_WIDTH-1:46*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_3_4_bottom;
			reg_valid_force_values[52*FORCE_EVAL_FIFO_DATA_WIDTH-1:51*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_1_mid;
			reg_valid_force_values[49*FORCE_EVAL_FIFO_DATA_WIDTH-1:48*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_1_top;
			reg_valid_force_values[51*FORCE_EVAL_FIFO_DATA_WIDTH-1:50*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_1_bottom;
			reg_valid_force_values[56*FORCE_EVAL_FIFO_DATA_WIDTH-1:55*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_2_mid;
			reg_valid_force_values[53*FORCE_EVAL_FIFO_DATA_WIDTH-1:52*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_2_top;
			reg_valid_force_values[55*FORCE_EVAL_FIFO_DATA_WIDTH-1:54*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_2_bottom;
			reg_valid_force_values[60*FORCE_EVAL_FIFO_DATA_WIDTH-1:59*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_3_mid;
			reg_valid_force_values[57*FORCE_EVAL_FIFO_DATA_WIDTH-1:56*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_3_top;
			reg_valid_force_values[59*FORCE_EVAL_FIFO_DATA_WIDTH-1:58*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_3_bottom;
			reg_valid_force_values[64*FORCE_EVAL_FIFO_DATA_WIDTH-1:63*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_4_mid;
			reg_valid_force_values[61*FORCE_EVAL_FIFO_DATA_WIDTH-1:60*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_4_top;
			reg_valid_force_values[63*FORCE_EVAL_FIFO_DATA_WIDTH-1:62*FORCE_EVAL_FIFO_DATA_WIDTH] = valid_force_values_4_4_bottom;
			end
		default:
			begin
			reg_valid_force_values = 0;
			end
	endcase
	end

always@(*)
	begin
	case(Arbitration_1_1_mid)
		6'b100000:
			begin
			valid_force_values_1_1_mid = ref_force_data_from_FIFO[1*FORCE_EVAL_FIFO_DATA_WIDTH-1:0*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b010000:
			begin
			valid_force_values_1_1_mid = neighbor_force_data_from_FIFO_1[1*FORCE_EVAL_FIFO_DATA_WIDTH-1:0*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_1_1_mid = neighbor_force_data_from_FIFO_1[4*FORCE_EVAL_FIFO_DATA_WIDTH-1:3*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_1_1_mid = neighbor_force_data_from_FIFO_1[14*FORCE_EVAL_FIFO_DATA_WIDTH-1:13*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_1_1_mid = neighbor_force_data_from_FIFO_2[13*FORCE_EVAL_FIFO_DATA_WIDTH-1:12*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_1_1_mid = neighbor_force_data_from_FIFO_2[16*FORCE_EVAL_FIFO_DATA_WIDTH-1:15*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_1_1_mid = 0;
			end
	endcase
	case(Arbitration_1_1_top)
		6'b100000:
			begin
			valid_force_values_1_1_top = 0;
			end
		6'b010000:
			begin
			valid_force_values_1_1_top = neighbor_force_data_from_FIFO_1[1*FORCE_EVAL_FIFO_DATA_WIDTH-1:0*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_1_1_top = neighbor_force_data_from_FIFO_1[4*FORCE_EVAL_FIFO_DATA_WIDTH-1:3*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_1_1_top = neighbor_force_data_from_FIFO_2[13*FORCE_EVAL_FIFO_DATA_WIDTH-1:12*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_1_1_top = neighbor_force_data_from_FIFO_2[14*FORCE_EVAL_FIFO_DATA_WIDTH-1:13*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_1_1_top = neighbor_force_data_from_FIFO_2[16*FORCE_EVAL_FIFO_DATA_WIDTH-1:15*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_1_1_top = 0;
			end
	endcase
	case(Arbitration_1_1_bottom)
		6'b100000:
			begin
			valid_force_values_1_1_bottom = 0;
			end
		6'b010000:
			begin
			valid_force_values_1_1_bottom = neighbor_force_data_from_FIFO_1[4*FORCE_EVAL_FIFO_DATA_WIDTH-1:3*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_1_1_bottom = neighbor_force_data_from_FIFO_1[14*FORCE_EVAL_FIFO_DATA_WIDTH-1:13*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_1_1_bottom = neighbor_force_data_from_FIFO_2[13*FORCE_EVAL_FIFO_DATA_WIDTH-1:12*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_1_1_bottom = neighbor_force_data_from_FIFO_2[16*FORCE_EVAL_FIFO_DATA_WIDTH-1:15*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_1_1_bottom = 0;
			end
		default:
			begin
			valid_force_values_1_1_bottom = 0;
			end
	endcase
	case(Arbitration_1_2_mid)
		6'b100000:
			begin
			valid_force_values_1_2_mid = ref_force_data_from_FIFO[2*FORCE_EVAL_FIFO_DATA_WIDTH-1:1*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b010000:
			begin
			valid_force_values_1_2_mid = neighbor_force_data_from_FIFO_1[1*FORCE_EVAL_FIFO_DATA_WIDTH-1:0*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_1_2_mid = neighbor_force_data_from_FIFO_1[2*FORCE_EVAL_FIFO_DATA_WIDTH-1:1*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_1_2_mid = neighbor_force_data_from_FIFO_1[15*FORCE_EVAL_FIFO_DATA_WIDTH-1:14*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_1_2_mid = neighbor_force_data_from_FIFO_2[13*FORCE_EVAL_FIFO_DATA_WIDTH-1:12*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_1_2_mid = neighbor_force_data_from_FIFO_2[14*FORCE_EVAL_FIFO_DATA_WIDTH-1:13*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_1_2_mid = 0;
			end
	endcase
	case(Arbitration_1_2_top)
		6'b100000:
			begin
			valid_force_values_1_2_top = 0;
			end
		6'b010000:
			begin
			valid_force_values_1_2_top = neighbor_force_data_from_FIFO_1[1*FORCE_EVAL_FIFO_DATA_WIDTH-1:0*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_1_2_top = neighbor_force_data_from_FIFO_1[2*FORCE_EVAL_FIFO_DATA_WIDTH-1:1*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_1_2_top = neighbor_force_data_from_FIFO_2[13*FORCE_EVAL_FIFO_DATA_WIDTH-1:12*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_1_2_top = neighbor_force_data_from_FIFO_2[14*FORCE_EVAL_FIFO_DATA_WIDTH-1:13*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_1_2_top = neighbor_force_data_from_FIFO_2[15*FORCE_EVAL_FIFO_DATA_WIDTH-1:14*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_1_2_top = 0;
			end
	endcase
	case(Arbitration_1_2_bottom)
		6'b100000:
			begin
			valid_force_values_1_2_bottom = 0;
			end
		6'b010000:
			begin
			valid_force_values_1_2_bottom = neighbor_force_data_from_FIFO_1[1*FORCE_EVAL_FIFO_DATA_WIDTH-1:0*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_1_2_bottom = neighbor_force_data_from_FIFO_1[15*FORCE_EVAL_FIFO_DATA_WIDTH-1:14*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_1_2_bottom = neighbor_force_data_from_FIFO_2[13*FORCE_EVAL_FIFO_DATA_WIDTH-1:12*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_1_2_bottom = neighbor_force_data_from_FIFO_2[14*FORCE_EVAL_FIFO_DATA_WIDTH-1:13*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_1_2_bottom = 0;
			end
		default:
			begin
			valid_force_values_1_2_bottom = 0;
			end
	endcase
	case(Arbitration_1_3_mid)
		6'b100000:
			begin
			valid_force_values_1_3_mid = ref_force_data_from_FIFO[3*FORCE_EVAL_FIFO_DATA_WIDTH-1:2*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b010000:
			begin
			valid_force_values_1_3_mid = neighbor_force_data_from_FIFO_1[2*FORCE_EVAL_FIFO_DATA_WIDTH-1:1*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_1_3_mid = neighbor_force_data_from_FIFO_1[3*FORCE_EVAL_FIFO_DATA_WIDTH-1:2*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_1_3_mid = neighbor_force_data_from_FIFO_1[16*FORCE_EVAL_FIFO_DATA_WIDTH-1:15*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_1_3_mid = neighbor_force_data_from_FIFO_2[14*FORCE_EVAL_FIFO_DATA_WIDTH-1:13*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_1_3_mid = neighbor_force_data_from_FIFO_2[15*FORCE_EVAL_FIFO_DATA_WIDTH-1:14*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_1_3_mid = 0;
			end
	endcase
	case(Arbitration_1_3_top)
		6'b100000:
			begin
			valid_force_values_1_3_top = 0;
			end
		6'b010000:
			begin
			valid_force_values_1_3_top = neighbor_force_data_from_FIFO_1[2*FORCE_EVAL_FIFO_DATA_WIDTH-1:1*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_1_3_top = neighbor_force_data_from_FIFO_1[3*FORCE_EVAL_FIFO_DATA_WIDTH-1:2*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_1_3_top = neighbor_force_data_from_FIFO_2[14*FORCE_EVAL_FIFO_DATA_WIDTH-1:13*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_1_3_top = neighbor_force_data_from_FIFO_2[15*FORCE_EVAL_FIFO_DATA_WIDTH-1:14*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_1_3_top = neighbor_force_data_from_FIFO_2[16*FORCE_EVAL_FIFO_DATA_WIDTH-1:15*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_1_3_top = 0;
			end
	endcase
	case(Arbitration_1_3_bottom)
		6'b100000:
			begin
			valid_force_values_1_3_bottom = 0;
			end
		6'b010000:
			begin
			valid_force_values_1_3_bottom = neighbor_force_data_from_FIFO_1[2*FORCE_EVAL_FIFO_DATA_WIDTH-1:1*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_1_3_bottom = neighbor_force_data_from_FIFO_1[16*FORCE_EVAL_FIFO_DATA_WIDTH-1:15*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_1_3_bottom = neighbor_force_data_from_FIFO_2[14*FORCE_EVAL_FIFO_DATA_WIDTH-1:13*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_1_3_bottom = neighbor_force_data_from_FIFO_2[15*FORCE_EVAL_FIFO_DATA_WIDTH-1:14*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_1_3_bottom = 0;
			end
		default:
			begin
			valid_force_values_1_3_bottom = 0;
			end
	endcase
	case(Arbitration_1_4_mid)
		6'b100000:
			begin
			valid_force_values_1_4_mid = ref_force_data_from_FIFO[4*FORCE_EVAL_FIFO_DATA_WIDTH-1:3*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b010000:
			begin
			valid_force_values_1_4_mid = neighbor_force_data_from_FIFO_1[3*FORCE_EVAL_FIFO_DATA_WIDTH-1:2*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_1_4_mid = neighbor_force_data_from_FIFO_1[4*FORCE_EVAL_FIFO_DATA_WIDTH-1:3*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_1_4_mid = neighbor_force_data_from_FIFO_1[13*FORCE_EVAL_FIFO_DATA_WIDTH-1:12*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_1_4_mid = neighbor_force_data_from_FIFO_2[15*FORCE_EVAL_FIFO_DATA_WIDTH-1:14*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_1_4_mid = neighbor_force_data_from_FIFO_2[16*FORCE_EVAL_FIFO_DATA_WIDTH-1:15*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_1_4_mid = 0;
			end
	endcase
	case(Arbitration_1_4_top)
		6'b100000:
			begin
			valid_force_values_1_4_top = 0;
			end
		6'b010000:
			begin
			valid_force_values_1_4_top = neighbor_force_data_from_FIFO_1[3*FORCE_EVAL_FIFO_DATA_WIDTH-1:2*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_1_4_top = neighbor_force_data_from_FIFO_1[4*FORCE_EVAL_FIFO_DATA_WIDTH-1:3*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_1_4_top = neighbor_force_data_from_FIFO_2[13*FORCE_EVAL_FIFO_DATA_WIDTH-1:12*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_1_4_top = neighbor_force_data_from_FIFO_2[15*FORCE_EVAL_FIFO_DATA_WIDTH-1:14*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_1_4_top = neighbor_force_data_from_FIFO_2[16*FORCE_EVAL_FIFO_DATA_WIDTH-1:15*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_1_4_top = 0;
			end
	endcase
	case(Arbitration_1_4_bottom)
		6'b100000:
			begin
			valid_force_values_1_4_bottom = 0;
			end
		6'b010000:
			begin
			valid_force_values_1_4_bottom = neighbor_force_data_from_FIFO_1[3*FORCE_EVAL_FIFO_DATA_WIDTH-1:2*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_1_4_bottom = neighbor_force_data_from_FIFO_1[13*FORCE_EVAL_FIFO_DATA_WIDTH-1:12*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_1_4_bottom = neighbor_force_data_from_FIFO_2[15*FORCE_EVAL_FIFO_DATA_WIDTH-1:14*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_1_4_bottom = neighbor_force_data_from_FIFO_2[16*FORCE_EVAL_FIFO_DATA_WIDTH-1:15*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_1_4_bottom = 0;
			end
		default:
			begin
			valid_force_values_1_4_bottom = 0;
			end
	endcase
	case(Arbitration_2_1_mid)
		6'b100000:
			begin
			valid_force_values_2_1_mid = ref_force_data_from_FIFO[5*FORCE_EVAL_FIFO_DATA_WIDTH-1:4*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b010000:
			begin
			valid_force_values_2_1_mid = neighbor_force_data_from_FIFO_1[2*FORCE_EVAL_FIFO_DATA_WIDTH-1:1*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_2_1_mid = neighbor_force_data_from_FIFO_1[5*FORCE_EVAL_FIFO_DATA_WIDTH-1:4*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_2_1_mid = neighbor_force_data_from_FIFO_1[8*FORCE_EVAL_FIFO_DATA_WIDTH-1:7*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_2_1_mid = neighbor_force_data_from_FIFO_2[1*FORCE_EVAL_FIFO_DATA_WIDTH-1:0*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_2_1_mid = neighbor_force_data_from_FIFO_2[4*FORCE_EVAL_FIFO_DATA_WIDTH-1:3*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_2_1_mid = 0;
			end
	endcase
	case(Arbitration_2_1_top)
		6'b100000:
			begin
			valid_force_values_2_1_top = 0;
			end
		6'b010000:
			begin
			valid_force_values_2_1_top = neighbor_force_data_from_FIFO_1[5*FORCE_EVAL_FIFO_DATA_WIDTH-1:4*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_2_1_top = neighbor_force_data_from_FIFO_1[8*FORCE_EVAL_FIFO_DATA_WIDTH-1:7*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_2_1_top = neighbor_force_data_from_FIFO_2[1*FORCE_EVAL_FIFO_DATA_WIDTH-1:0*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_2_1_top = neighbor_force_data_from_FIFO_2[2*FORCE_EVAL_FIFO_DATA_WIDTH-1:1*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_2_1_top = neighbor_force_data_from_FIFO_2[4*FORCE_EVAL_FIFO_DATA_WIDTH-1:3*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_2_1_top = 0;
			end
	endcase
	case(Arbitration_2_1_bottom)
		6'b100000:
			begin
			valid_force_values_2_1_bottom = 0;
			end
		6'b010000:
			begin
			valid_force_values_2_1_bottom = neighbor_force_data_from_FIFO_1[2*FORCE_EVAL_FIFO_DATA_WIDTH-1:1*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_2_1_bottom = neighbor_force_data_from_FIFO_1[8*FORCE_EVAL_FIFO_DATA_WIDTH-1:7*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_2_1_bottom = neighbor_force_data_from_FIFO_2[1*FORCE_EVAL_FIFO_DATA_WIDTH-1:0*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_2_1_bottom = neighbor_force_data_from_FIFO_2[4*FORCE_EVAL_FIFO_DATA_WIDTH-1:3*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_2_1_bottom = 0;
			end
		default:
			begin
			valid_force_values_2_1_bottom = 0;
			end
	endcase
	case(Arbitration_2_2_mid)
		6'b100000:
			begin
			valid_force_values_2_2_mid = ref_force_data_from_FIFO[6*FORCE_EVAL_FIFO_DATA_WIDTH-1:5*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b010000:
			begin
			valid_force_values_2_2_mid = neighbor_force_data_from_FIFO_1[3*FORCE_EVAL_FIFO_DATA_WIDTH-1:2*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_2_2_mid = neighbor_force_data_from_FIFO_1[5*FORCE_EVAL_FIFO_DATA_WIDTH-1:4*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_2_2_mid = neighbor_force_data_from_FIFO_1[6*FORCE_EVAL_FIFO_DATA_WIDTH-1:5*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_2_2_mid = neighbor_force_data_from_FIFO_2[1*FORCE_EVAL_FIFO_DATA_WIDTH-1:0*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_2_2_mid = neighbor_force_data_from_FIFO_2[2*FORCE_EVAL_FIFO_DATA_WIDTH-1:1*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_2_2_mid = 0;
			end
	endcase
	case(Arbitration_2_2_top)
		6'b100000:
			begin
			valid_force_values_2_2_top = 0;
			end
		6'b010000:
			begin
			valid_force_values_2_2_top = neighbor_force_data_from_FIFO_1[5*FORCE_EVAL_FIFO_DATA_WIDTH-1:4*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_2_2_top = neighbor_force_data_from_FIFO_1[6*FORCE_EVAL_FIFO_DATA_WIDTH-1:5*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_2_2_top = neighbor_force_data_from_FIFO_2[1*FORCE_EVAL_FIFO_DATA_WIDTH-1:0*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_2_2_top = neighbor_force_data_from_FIFO_2[2*FORCE_EVAL_FIFO_DATA_WIDTH-1:1*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_2_2_top = neighbor_force_data_from_FIFO_2[3*FORCE_EVAL_FIFO_DATA_WIDTH-1:2*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_2_2_top = 0;
			end
	endcase
	case(Arbitration_2_2_bottom)
		6'b100000:
			begin
			valid_force_values_2_2_bottom = 0;
			end
		6'b010000:
			begin
			valid_force_values_2_2_bottom = neighbor_force_data_from_FIFO_1[3*FORCE_EVAL_FIFO_DATA_WIDTH-1:2*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_2_2_bottom = neighbor_force_data_from_FIFO_1[5*FORCE_EVAL_FIFO_DATA_WIDTH-1:4*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_2_2_bottom = neighbor_force_data_from_FIFO_2[1*FORCE_EVAL_FIFO_DATA_WIDTH-1:0*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_2_2_bottom = neighbor_force_data_from_FIFO_2[2*FORCE_EVAL_FIFO_DATA_WIDTH-1:1*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_2_2_bottom = 0;
			end
		default:
			begin
			valid_force_values_2_2_bottom = 0;
			end
	endcase
	case(Arbitration_2_3_mid)
		6'b100000:
			begin
			valid_force_values_2_3_mid = ref_force_data_from_FIFO[7*FORCE_EVAL_FIFO_DATA_WIDTH-1:6*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b010000:
			begin
			valid_force_values_2_3_mid = neighbor_force_data_from_FIFO_1[4*FORCE_EVAL_FIFO_DATA_WIDTH-1:3*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_2_3_mid = neighbor_force_data_from_FIFO_1[6*FORCE_EVAL_FIFO_DATA_WIDTH-1:5*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_2_3_mid = neighbor_force_data_from_FIFO_1[7*FORCE_EVAL_FIFO_DATA_WIDTH-1:6*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_2_3_mid = neighbor_force_data_from_FIFO_2[2*FORCE_EVAL_FIFO_DATA_WIDTH-1:1*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_2_3_mid = neighbor_force_data_from_FIFO_2[3*FORCE_EVAL_FIFO_DATA_WIDTH-1:2*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_2_3_mid = 0;
			end
	endcase
	case(Arbitration_2_3_top)
		6'b100000:
			begin
			valid_force_values_2_3_top = 0;
			end
		6'b010000:
			begin
			valid_force_values_2_3_top = neighbor_force_data_from_FIFO_1[6*FORCE_EVAL_FIFO_DATA_WIDTH-1:5*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_2_3_top = neighbor_force_data_from_FIFO_1[7*FORCE_EVAL_FIFO_DATA_WIDTH-1:6*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_2_3_top = neighbor_force_data_from_FIFO_2[2*FORCE_EVAL_FIFO_DATA_WIDTH-1:1*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_2_3_top = neighbor_force_data_from_FIFO_2[3*FORCE_EVAL_FIFO_DATA_WIDTH-1:2*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_2_3_top = neighbor_force_data_from_FIFO_2[4*FORCE_EVAL_FIFO_DATA_WIDTH-1:3*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_2_3_top = 0;
			end
	endcase
	case(Arbitration_2_3_bottom)
		6'b100000:
			begin
			valid_force_values_2_3_bottom = 0;
			end
		6'b010000:
			begin
			valid_force_values_2_3_bottom = neighbor_force_data_from_FIFO_1[4*FORCE_EVAL_FIFO_DATA_WIDTH-1:3*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_2_3_bottom = neighbor_force_data_from_FIFO_1[6*FORCE_EVAL_FIFO_DATA_WIDTH-1:5*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_2_3_bottom = neighbor_force_data_from_FIFO_2[2*FORCE_EVAL_FIFO_DATA_WIDTH-1:1*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_2_3_bottom = neighbor_force_data_from_FIFO_2[3*FORCE_EVAL_FIFO_DATA_WIDTH-1:2*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_2_3_bottom = 0;
			end
		default:
			begin
			valid_force_values_2_3_bottom = 0;
			end
	endcase
	case(Arbitration_2_4_mid)
		6'b100000:
			begin
			valid_force_values_2_4_mid = ref_force_data_from_FIFO[8*FORCE_EVAL_FIFO_DATA_WIDTH-1:7*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b010000:
			begin
			valid_force_values_2_4_mid = neighbor_force_data_from_FIFO_1[1*FORCE_EVAL_FIFO_DATA_WIDTH-1:0*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_2_4_mid = neighbor_force_data_from_FIFO_1[7*FORCE_EVAL_FIFO_DATA_WIDTH-1:6*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_2_4_mid = neighbor_force_data_from_FIFO_1[8*FORCE_EVAL_FIFO_DATA_WIDTH-1:7*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_2_4_mid = neighbor_force_data_from_FIFO_2[3*FORCE_EVAL_FIFO_DATA_WIDTH-1:2*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_2_4_mid = neighbor_force_data_from_FIFO_2[4*FORCE_EVAL_FIFO_DATA_WIDTH-1:3*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_2_4_mid = 0;
			end
	endcase
	case(Arbitration_2_4_top)
		6'b100000:
			begin
			valid_force_values_2_4_top = 0;
			end
		6'b010000:
			begin
			valid_force_values_2_4_top = neighbor_force_data_from_FIFO_1[7*FORCE_EVAL_FIFO_DATA_WIDTH-1:6*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_2_4_top = neighbor_force_data_from_FIFO_1[8*FORCE_EVAL_FIFO_DATA_WIDTH-1:7*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_2_4_top = neighbor_force_data_from_FIFO_2[1*FORCE_EVAL_FIFO_DATA_WIDTH-1:0*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_2_4_top = neighbor_force_data_from_FIFO_2[3*FORCE_EVAL_FIFO_DATA_WIDTH-1:2*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_2_4_top = neighbor_force_data_from_FIFO_2[4*FORCE_EVAL_FIFO_DATA_WIDTH-1:3*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_2_4_top = 0;
			end
	endcase
	case(Arbitration_2_4_bottom)
		6'b100000:
			begin
			valid_force_values_2_4_bottom = 0;
			end
		6'b010000:
			begin
			valid_force_values_2_4_bottom = neighbor_force_data_from_FIFO_1[1*FORCE_EVAL_FIFO_DATA_WIDTH-1:0*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_2_4_bottom = neighbor_force_data_from_FIFO_1[7*FORCE_EVAL_FIFO_DATA_WIDTH-1:6*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_2_4_bottom = neighbor_force_data_from_FIFO_2[3*FORCE_EVAL_FIFO_DATA_WIDTH-1:2*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_2_4_bottom = neighbor_force_data_from_FIFO_2[4*FORCE_EVAL_FIFO_DATA_WIDTH-1:3*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_2_4_bottom = 0;
			end
		default:
			begin
			valid_force_values_2_4_bottom = 0;
			end
	endcase
	case(Arbitration_3_1_mid)
		6'b100000:
			begin
			valid_force_values_3_1_mid = ref_force_data_from_FIFO[9*FORCE_EVAL_FIFO_DATA_WIDTH-1:8*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b010000:
			begin
			valid_force_values_3_1_mid = neighbor_force_data_from_FIFO_1[6*FORCE_EVAL_FIFO_DATA_WIDTH-1:5*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_3_1_mid = neighbor_force_data_from_FIFO_1[9*FORCE_EVAL_FIFO_DATA_WIDTH-1:8*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_3_1_mid = neighbor_force_data_from_FIFO_1[12*FORCE_EVAL_FIFO_DATA_WIDTH-1:11*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_3_1_mid = neighbor_force_data_from_FIFO_2[5*FORCE_EVAL_FIFO_DATA_WIDTH-1:4*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_3_1_mid = neighbor_force_data_from_FIFO_2[8*FORCE_EVAL_FIFO_DATA_WIDTH-1:7*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_3_1_mid = 0;
			end
	endcase
	case(Arbitration_3_1_top)
		6'b100000:
			begin
			valid_force_values_3_1_top = 0;
			end
		6'b010000:
			begin
			valid_force_values_3_1_top = neighbor_force_data_from_FIFO_1[9*FORCE_EVAL_FIFO_DATA_WIDTH-1:8*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_3_1_top = neighbor_force_data_from_FIFO_1[12*FORCE_EVAL_FIFO_DATA_WIDTH-1:11*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_3_1_top = neighbor_force_data_from_FIFO_2[5*FORCE_EVAL_FIFO_DATA_WIDTH-1:4*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_3_1_top = neighbor_force_data_from_FIFO_2[6*FORCE_EVAL_FIFO_DATA_WIDTH-1:5*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_3_1_top = neighbor_force_data_from_FIFO_2[8*FORCE_EVAL_FIFO_DATA_WIDTH-1:7*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_3_1_top = 0;
			end
	endcase
	case(Arbitration_3_1_bottom)
		6'b100000:
			begin
			valid_force_values_3_1_bottom = 0;
			end
		6'b010000:
			begin
			valid_force_values_3_1_bottom = neighbor_force_data_from_FIFO_1[6*FORCE_EVAL_FIFO_DATA_WIDTH-1:5*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_3_1_bottom = neighbor_force_data_from_FIFO_1[12*FORCE_EVAL_FIFO_DATA_WIDTH-1:11*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_3_1_bottom = neighbor_force_data_from_FIFO_2[5*FORCE_EVAL_FIFO_DATA_WIDTH-1:4*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_3_1_bottom = neighbor_force_data_from_FIFO_2[8*FORCE_EVAL_FIFO_DATA_WIDTH-1:7*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_3_1_bottom = 0;
			end
		default:
			begin
			valid_force_values_3_1_bottom = 0;
			end
	endcase
	case(Arbitration_3_2_mid)
		6'b100000:
			begin
			valid_force_values_3_2_mid = ref_force_data_from_FIFO[10*FORCE_EVAL_FIFO_DATA_WIDTH-1:9*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b010000:
			begin
			valid_force_values_3_2_mid = neighbor_force_data_from_FIFO_1[7*FORCE_EVAL_FIFO_DATA_WIDTH-1:6*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_3_2_mid = neighbor_force_data_from_FIFO_1[9*FORCE_EVAL_FIFO_DATA_WIDTH-1:8*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_3_2_mid = neighbor_force_data_from_FIFO_1[10*FORCE_EVAL_FIFO_DATA_WIDTH-1:9*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_3_2_mid = neighbor_force_data_from_FIFO_2[5*FORCE_EVAL_FIFO_DATA_WIDTH-1:4*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_3_2_mid = neighbor_force_data_from_FIFO_2[6*FORCE_EVAL_FIFO_DATA_WIDTH-1:5*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_3_2_mid = 0;
			end
	endcase
	case(Arbitration_3_2_top)
		6'b100000:
			begin
			valid_force_values_3_2_top = 0;
			end
		6'b010000:
			begin
			valid_force_values_3_2_top = neighbor_force_data_from_FIFO_1[9*FORCE_EVAL_FIFO_DATA_WIDTH-1:8*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_3_2_top = neighbor_force_data_from_FIFO_1[10*FORCE_EVAL_FIFO_DATA_WIDTH-1:9*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_3_2_top = neighbor_force_data_from_FIFO_2[5*FORCE_EVAL_FIFO_DATA_WIDTH-1:4*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_3_2_top = neighbor_force_data_from_FIFO_2[6*FORCE_EVAL_FIFO_DATA_WIDTH-1:5*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_3_2_top = neighbor_force_data_from_FIFO_2[7*FORCE_EVAL_FIFO_DATA_WIDTH-1:6*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_3_2_top = 0;
			end
	endcase
	case(Arbitration_3_2_bottom)
		6'b100000:
			begin
			valid_force_values_3_2_bottom = 0;
			end
		6'b010000:
			begin
			valid_force_values_3_2_bottom = neighbor_force_data_from_FIFO_1[7*FORCE_EVAL_FIFO_DATA_WIDTH-1:6*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_3_2_bottom = neighbor_force_data_from_FIFO_1[9*FORCE_EVAL_FIFO_DATA_WIDTH-1:8*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_3_2_bottom = neighbor_force_data_from_FIFO_2[5*FORCE_EVAL_FIFO_DATA_WIDTH-1:4*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_3_2_bottom = neighbor_force_data_from_FIFO_2[6*FORCE_EVAL_FIFO_DATA_WIDTH-1:5*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_3_2_bottom = 0;
			end
		default:
			begin
			valid_force_values_3_2_bottom = 0;
			end
	endcase
	case(Arbitration_3_3_mid)
		6'b100000:
			begin
			valid_force_values_3_3_mid = ref_force_data_from_FIFO[11*FORCE_EVAL_FIFO_DATA_WIDTH-1:10*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b010000:
			begin
			valid_force_values_3_3_mid = neighbor_force_data_from_FIFO_1[8*FORCE_EVAL_FIFO_DATA_WIDTH-1:7*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_3_3_mid = neighbor_force_data_from_FIFO_1[10*FORCE_EVAL_FIFO_DATA_WIDTH-1:9*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_3_3_mid = neighbor_force_data_from_FIFO_1[11*FORCE_EVAL_FIFO_DATA_WIDTH-1:10*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_3_3_mid = neighbor_force_data_from_FIFO_2[6*FORCE_EVAL_FIFO_DATA_WIDTH-1:5*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_3_3_mid = neighbor_force_data_from_FIFO_2[7*FORCE_EVAL_FIFO_DATA_WIDTH-1:6*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_3_3_mid = 0;
			end
	endcase
	case(Arbitration_3_3_top)
		6'b100000:
			begin
			valid_force_values_3_3_top = 0;
			end
		6'b010000:
			begin
			valid_force_values_3_3_top = neighbor_force_data_from_FIFO_1[10*FORCE_EVAL_FIFO_DATA_WIDTH-1:9*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_3_3_top = neighbor_force_data_from_FIFO_1[11*FORCE_EVAL_FIFO_DATA_WIDTH-1:10*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_3_3_top = neighbor_force_data_from_FIFO_2[6*FORCE_EVAL_FIFO_DATA_WIDTH-1:5*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_3_3_top = neighbor_force_data_from_FIFO_2[7*FORCE_EVAL_FIFO_DATA_WIDTH-1:6*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_3_3_top = neighbor_force_data_from_FIFO_2[8*FORCE_EVAL_FIFO_DATA_WIDTH-1:7*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_3_3_top = 0;
			end
	endcase
	case(Arbitration_3_3_bottom)
		6'b100000:
			begin
			valid_force_values_3_3_bottom = 0;
			end
		6'b010000:
			begin
			valid_force_values_3_3_bottom = neighbor_force_data_from_FIFO_1[8*FORCE_EVAL_FIFO_DATA_WIDTH-1:7*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_3_3_bottom = neighbor_force_data_from_FIFO_1[10*FORCE_EVAL_FIFO_DATA_WIDTH-1:9*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_3_3_bottom = neighbor_force_data_from_FIFO_2[6*FORCE_EVAL_FIFO_DATA_WIDTH-1:5*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_3_3_bottom = neighbor_force_data_from_FIFO_2[7*FORCE_EVAL_FIFO_DATA_WIDTH-1:6*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_3_3_bottom = 0;
			end
		default:
			begin
			valid_force_values_3_3_bottom = 0;
			end
	endcase
	case(Arbitration_3_4_mid)
		6'b100000:
			begin
			valid_force_values_3_4_mid = ref_force_data_from_FIFO[12*FORCE_EVAL_FIFO_DATA_WIDTH-1:11*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b010000:
			begin
			valid_force_values_3_4_mid = neighbor_force_data_from_FIFO_1[5*FORCE_EVAL_FIFO_DATA_WIDTH-1:4*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_3_4_mid = neighbor_force_data_from_FIFO_1[11*FORCE_EVAL_FIFO_DATA_WIDTH-1:10*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_3_4_mid = neighbor_force_data_from_FIFO_1[12*FORCE_EVAL_FIFO_DATA_WIDTH-1:11*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_3_4_mid = neighbor_force_data_from_FIFO_2[7*FORCE_EVAL_FIFO_DATA_WIDTH-1:6*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_3_4_mid = neighbor_force_data_from_FIFO_2[8*FORCE_EVAL_FIFO_DATA_WIDTH-1:7*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_3_4_mid = 0;
			end
	endcase
	case(Arbitration_3_4_top)
		6'b100000:
			begin
			valid_force_values_3_4_top = 0;
			end
		6'b010000:
			begin
			valid_force_values_3_4_top = neighbor_force_data_from_FIFO_1[11*FORCE_EVAL_FIFO_DATA_WIDTH-1:10*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_3_4_top = neighbor_force_data_from_FIFO_1[12*FORCE_EVAL_FIFO_DATA_WIDTH-1:11*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_3_4_top = neighbor_force_data_from_FIFO_2[5*FORCE_EVAL_FIFO_DATA_WIDTH-1:4*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_3_4_top = neighbor_force_data_from_FIFO_2[7*FORCE_EVAL_FIFO_DATA_WIDTH-1:6*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_3_4_top = neighbor_force_data_from_FIFO_2[8*FORCE_EVAL_FIFO_DATA_WIDTH-1:7*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_3_4_top = 0;
			end
	endcase
	case(Arbitration_3_4_bottom)
		6'b100000:
			begin
			valid_force_values_3_4_bottom = 0;
			end
		6'b010000:
			begin
			valid_force_values_3_4_bottom = neighbor_force_data_from_FIFO_1[5*FORCE_EVAL_FIFO_DATA_WIDTH-1:4*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_3_4_bottom = neighbor_force_data_from_FIFO_1[11*FORCE_EVAL_FIFO_DATA_WIDTH-1:10*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_3_4_bottom = neighbor_force_data_from_FIFO_2[7*FORCE_EVAL_FIFO_DATA_WIDTH-1:6*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_3_4_bottom = neighbor_force_data_from_FIFO_2[8*FORCE_EVAL_FIFO_DATA_WIDTH-1:7*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_3_4_bottom = 0;
			end
		default:
			begin
			valid_force_values_3_4_bottom = 0;
			end
	endcase
	case(Arbitration_4_1_mid)
		6'b100000:
			begin
			valid_force_values_4_1_mid = ref_force_data_from_FIFO[13*FORCE_EVAL_FIFO_DATA_WIDTH-1:12*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b010000:
			begin
			valid_force_values_4_1_mid = neighbor_force_data_from_FIFO_1[10*FORCE_EVAL_FIFO_DATA_WIDTH-1:9*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_4_1_mid = neighbor_force_data_from_FIFO_1[13*FORCE_EVAL_FIFO_DATA_WIDTH-1:12*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_4_1_mid = neighbor_force_data_from_FIFO_1[16*FORCE_EVAL_FIFO_DATA_WIDTH-1:15*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_4_1_mid = neighbor_force_data_from_FIFO_2[9*FORCE_EVAL_FIFO_DATA_WIDTH-1:8*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_4_1_mid = neighbor_force_data_from_FIFO_2[12*FORCE_EVAL_FIFO_DATA_WIDTH-1:11*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_4_1_mid = 0;
			end
	endcase
	case(Arbitration_4_1_top)
		6'b100000:
			begin
			valid_force_values_4_1_top = 0;
			end
		6'b010000:
			begin
			valid_force_values_4_1_top = neighbor_force_data_from_FIFO_1[13*FORCE_EVAL_FIFO_DATA_WIDTH-1:12*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_4_1_top = neighbor_force_data_from_FIFO_1[16*FORCE_EVAL_FIFO_DATA_WIDTH-1:15*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_4_1_top = neighbor_force_data_from_FIFO_2[9*FORCE_EVAL_FIFO_DATA_WIDTH-1:8*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_4_1_top = neighbor_force_data_from_FIFO_2[10*FORCE_EVAL_FIFO_DATA_WIDTH-1:9*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_4_1_top = neighbor_force_data_from_FIFO_2[12*FORCE_EVAL_FIFO_DATA_WIDTH-1:11*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_4_1_top = 0;
			end
	endcase
	case(Arbitration_4_1_bottom)
		6'b100000:
			begin
			valid_force_values_4_1_bottom = 0;
			end
		6'b010000:
			begin
			valid_force_values_4_1_bottom = neighbor_force_data_from_FIFO_1[10*FORCE_EVAL_FIFO_DATA_WIDTH-1:9*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_4_1_bottom = neighbor_force_data_from_FIFO_1[16*FORCE_EVAL_FIFO_DATA_WIDTH-1:15*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_4_1_bottom = neighbor_force_data_from_FIFO_2[9*FORCE_EVAL_FIFO_DATA_WIDTH-1:8*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_4_1_bottom = neighbor_force_data_from_FIFO_2[12*FORCE_EVAL_FIFO_DATA_WIDTH-1:11*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_4_1_bottom = 0;
			end
		default:
			begin
			valid_force_values_4_1_bottom = 0;
			end
	endcase
	case(Arbitration_4_2_mid)
		6'b100000:
			begin
			valid_force_values_4_2_mid = ref_force_data_from_FIFO[14*FORCE_EVAL_FIFO_DATA_WIDTH-1:13*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b010000:
			begin
			valid_force_values_4_2_mid = neighbor_force_data_from_FIFO_1[11*FORCE_EVAL_FIFO_DATA_WIDTH-1:10*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_4_2_mid = neighbor_force_data_from_FIFO_1[13*FORCE_EVAL_FIFO_DATA_WIDTH-1:12*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_4_2_mid = neighbor_force_data_from_FIFO_1[14*FORCE_EVAL_FIFO_DATA_WIDTH-1:13*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_4_2_mid = neighbor_force_data_from_FIFO_2[9*FORCE_EVAL_FIFO_DATA_WIDTH-1:8*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_4_2_mid = neighbor_force_data_from_FIFO_2[10*FORCE_EVAL_FIFO_DATA_WIDTH-1:9*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_4_2_mid = 0;
			end
	endcase
	case(Arbitration_4_2_top)
		6'b100000:
			begin
			valid_force_values_4_2_top = 0;
			end
		6'b010000:
			begin
			valid_force_values_4_2_top = neighbor_force_data_from_FIFO_1[13*FORCE_EVAL_FIFO_DATA_WIDTH-1:12*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_4_2_top = neighbor_force_data_from_FIFO_1[14*FORCE_EVAL_FIFO_DATA_WIDTH-1:13*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_4_2_top = neighbor_force_data_from_FIFO_2[9*FORCE_EVAL_FIFO_DATA_WIDTH-1:8*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_4_2_top = neighbor_force_data_from_FIFO_2[10*FORCE_EVAL_FIFO_DATA_WIDTH-1:9*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_4_2_top = neighbor_force_data_from_FIFO_2[11*FORCE_EVAL_FIFO_DATA_WIDTH-1:10*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_4_2_top = 0;
			end
	endcase
	case(Arbitration_4_2_bottom)
		6'b100000:
			begin
			valid_force_values_4_2_bottom = 0;
			end
		6'b010000:
			begin
			valid_force_values_4_2_bottom = neighbor_force_data_from_FIFO_1[11*FORCE_EVAL_FIFO_DATA_WIDTH-1:10*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_4_2_bottom = neighbor_force_data_from_FIFO_1[13*FORCE_EVAL_FIFO_DATA_WIDTH-1:12*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_4_2_bottom = neighbor_force_data_from_FIFO_2[9*FORCE_EVAL_FIFO_DATA_WIDTH-1:8*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_4_2_bottom = neighbor_force_data_from_FIFO_2[10*FORCE_EVAL_FIFO_DATA_WIDTH-1:9*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_4_2_bottom = 0;
			end
		default:
			begin
			valid_force_values_4_2_bottom = 0;
			end
	endcase
	case(Arbitration_4_3_mid)
		6'b100000:
			begin
			valid_force_values_4_3_mid = ref_force_data_from_FIFO[15*FORCE_EVAL_FIFO_DATA_WIDTH-1:14*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b010000:
			begin
			valid_force_values_4_3_mid = neighbor_force_data_from_FIFO_1[12*FORCE_EVAL_FIFO_DATA_WIDTH-1:11*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_4_3_mid = neighbor_force_data_from_FIFO_1[14*FORCE_EVAL_FIFO_DATA_WIDTH-1:13*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_4_3_mid = neighbor_force_data_from_FIFO_1[15*FORCE_EVAL_FIFO_DATA_WIDTH-1:14*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_4_3_mid = neighbor_force_data_from_FIFO_2[10*FORCE_EVAL_FIFO_DATA_WIDTH-1:9*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_4_3_mid = neighbor_force_data_from_FIFO_2[11*FORCE_EVAL_FIFO_DATA_WIDTH-1:10*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_4_3_mid = 0;
			end
	endcase
	case(Arbitration_4_3_top)
		6'b100000:
			begin
			valid_force_values_4_3_top = 0;
			end
		6'b010000:
			begin
			valid_force_values_4_3_top = neighbor_force_data_from_FIFO_1[14*FORCE_EVAL_FIFO_DATA_WIDTH-1:13*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_4_3_top = neighbor_force_data_from_FIFO_1[15*FORCE_EVAL_FIFO_DATA_WIDTH-1:14*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_4_3_top = neighbor_force_data_from_FIFO_2[10*FORCE_EVAL_FIFO_DATA_WIDTH-1:9*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_4_3_top = neighbor_force_data_from_FIFO_2[11*FORCE_EVAL_FIFO_DATA_WIDTH-1:10*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_4_3_top = neighbor_force_data_from_FIFO_2[12*FORCE_EVAL_FIFO_DATA_WIDTH-1:11*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_4_3_top = 0;
			end
	endcase
	case(Arbitration_4_3_bottom)
		6'b100000:
			begin
			valid_force_values_4_3_bottom = 0;
			end
		6'b010000:
			begin
			valid_force_values_4_3_bottom = neighbor_force_data_from_FIFO_1[12*FORCE_EVAL_FIFO_DATA_WIDTH-1:11*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_4_3_bottom = neighbor_force_data_from_FIFO_1[14*FORCE_EVAL_FIFO_DATA_WIDTH-1:13*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_4_3_bottom = neighbor_force_data_from_FIFO_2[10*FORCE_EVAL_FIFO_DATA_WIDTH-1:9*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_4_3_bottom = neighbor_force_data_from_FIFO_2[11*FORCE_EVAL_FIFO_DATA_WIDTH-1:10*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_4_3_bottom = 0;
			end
		default:
			begin
			valid_force_values_4_3_bottom = 0;
			end
	endcase
	case(Arbitration_4_4_mid)
		6'b100000:
			begin
			valid_force_values_4_4_mid = ref_force_data_from_FIFO[16*FORCE_EVAL_FIFO_DATA_WIDTH-1:15*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b010000:
			begin
			valid_force_values_4_4_mid = neighbor_force_data_from_FIFO_1[9*FORCE_EVAL_FIFO_DATA_WIDTH-1:8*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_4_4_mid = neighbor_force_data_from_FIFO_1[15*FORCE_EVAL_FIFO_DATA_WIDTH-1:14*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_4_4_mid = neighbor_force_data_from_FIFO_1[16*FORCE_EVAL_FIFO_DATA_WIDTH-1:15*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_4_4_mid = neighbor_force_data_from_FIFO_2[11*FORCE_EVAL_FIFO_DATA_WIDTH-1:10*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_4_4_mid = neighbor_force_data_from_FIFO_2[12*FORCE_EVAL_FIFO_DATA_WIDTH-1:11*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_4_4_mid = 0;
			end
	endcase
	case(Arbitration_4_4_top)
		6'b100000:
			begin
			valid_force_values_4_4_top = 0;
			end
		6'b010000:
			begin
			valid_force_values_4_4_top = neighbor_force_data_from_FIFO_1[15*FORCE_EVAL_FIFO_DATA_WIDTH-1:14*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_4_4_top = neighbor_force_data_from_FIFO_1[16*FORCE_EVAL_FIFO_DATA_WIDTH-1:15*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_4_4_top = neighbor_force_data_from_FIFO_2[9*FORCE_EVAL_FIFO_DATA_WIDTH-1:8*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_4_4_top = neighbor_force_data_from_FIFO_2[11*FORCE_EVAL_FIFO_DATA_WIDTH-1:10*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_4_4_top = neighbor_force_data_from_FIFO_2[12*FORCE_EVAL_FIFO_DATA_WIDTH-1:11*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		default:
			begin
			valid_force_values_4_4_top = 0;
			end
	endcase
	case(Arbitration_4_4_bottom)
		6'b100000:
			begin
			valid_force_values_4_4_bottom = 0;
			end
		6'b010000:
			begin
			valid_force_values_4_4_bottom = neighbor_force_data_from_FIFO_1[9*FORCE_EVAL_FIFO_DATA_WIDTH-1:8*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b001000:
			begin
			valid_force_values_4_4_bottom = neighbor_force_data_from_FIFO_1[15*FORCE_EVAL_FIFO_DATA_WIDTH-1:14*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000100:
			begin
			valid_force_values_4_4_bottom = neighbor_force_data_from_FIFO_2[11*FORCE_EVAL_FIFO_DATA_WIDTH-1:10*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000010:
			begin
			valid_force_values_4_4_bottom = neighbor_force_data_from_FIFO_2[12*FORCE_EVAL_FIFO_DATA_WIDTH-1:11*FORCE_EVAL_FIFO_DATA_WIDTH];
			end
		6'b000001:
			begin
			valid_force_values_4_4_bottom = 0;
			end
		default:
			begin
			valid_force_values_4_4_bottom = 0;
			end
	endcase
	end

always@(*)
	begin
	case(neighbor_force_data_from_FIFO_1[0*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:0*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_222:
			begin
			force_valid_1_1_mid_1 = neighbor_force_valid_1[0];
			force_valid_1_1_top_1 = 1'b0;
			force_valid_1_2_bottom_1 = 1'b0;
			force_valid_1_2_mid_1 = 1'b0;
			force_valid_1_2_top_1 = 1'b0;
			force_valid_2_4_bottom_1 = 1'b0;
			force_valid_2_4_mid_1 = 1'b0;
			end
		BINARY_223:
			begin
			force_valid_1_1_top_1 = neighbor_force_valid_1[0];
			force_valid_1_1_mid_1 = 1'b0;
			force_valid_1_2_bottom_1 = 1'b0;
			force_valid_1_2_mid_1 = 1'b0;
			force_valid_1_2_top_1 = 1'b0;
			force_valid_2_4_bottom_1 = 1'b0;
			force_valid_2_4_mid_1 = 1'b0;
			end
		BINARY_231:
			begin
			force_valid_1_2_bottom_1 = neighbor_force_valid_1[0];
			force_valid_1_1_mid_1 = 1'b0;
			force_valid_1_1_top_1 = 1'b0;
			force_valid_1_2_mid_1 = 1'b0;
			force_valid_1_2_top_1 = 1'b0;
			force_valid_2_4_bottom_1 = 1'b0;
			force_valid_2_4_mid_1 = 1'b0;
			end
		BINARY_232:
			begin
			force_valid_1_2_mid_1 = neighbor_force_valid_1[0];
			force_valid_1_1_mid_1 = 1'b0;
			force_valid_1_1_top_1 = 1'b0;
			force_valid_1_2_bottom_1 = 1'b0;
			force_valid_1_2_top_1 = 1'b0;
			force_valid_2_4_bottom_1 = 1'b0;
			force_valid_2_4_mid_1 = 1'b0;
			end
		BINARY_233:
			begin
			force_valid_1_2_top_1 = neighbor_force_valid_1[0];
			force_valid_1_1_mid_1 = 1'b0;
			force_valid_1_1_top_1 = 1'b0;
			force_valid_1_2_bottom_1 = 1'b0;
			force_valid_1_2_mid_1 = 1'b0;
			force_valid_2_4_bottom_1 = 1'b0;
			force_valid_2_4_mid_1 = 1'b0;
			end
		BINARY_311:
			begin
			force_valid_2_4_bottom_1 = neighbor_force_valid_1[0];
			force_valid_1_1_mid_1 = 1'b0;
			force_valid_1_1_top_1 = 1'b0;
			force_valid_1_2_bottom_1 = 1'b0;
			force_valid_1_2_mid_1 = 1'b0;
			force_valid_1_2_top_1 = 1'b0;
			force_valid_2_4_mid_1 = 1'b0;
			end
		BINARY_312:
			begin
			force_valid_2_4_mid_1 = neighbor_force_valid_1[0];
			force_valid_1_1_mid_1 = 1'b0;
			force_valid_1_1_top_1 = 1'b0;
			force_valid_1_2_bottom_1 = 1'b0;
			force_valid_1_2_mid_1 = 1'b0;
			force_valid_1_2_top_1 = 1'b0;
			force_valid_2_4_bottom_1 = 1'b0;
			end
		default:
			begin
			force_valid_1_1_mid_1 = 1'b0;
			force_valid_1_1_top_1 = 1'b0;
			force_valid_1_2_bottom_1 = 1'b0;
			force_valid_1_2_mid_1 = 1'b0;
			force_valid_1_2_top_1 = 1'b0;
			force_valid_2_4_bottom_1 = 1'b0;
			force_valid_2_4_mid_1 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_1[1*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:1*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_222:
			begin
			force_valid_1_2_mid_2 = neighbor_force_valid_1[1];
			force_valid_1_2_top_2 = 1'b0;
			force_valid_1_3_bottom_1 = 1'b0;
			force_valid_1_3_mid_1 = 1'b0;
			force_valid_1_3_top_1 = 1'b0;
			force_valid_2_1_bottom_1 = 1'b0;
			force_valid_2_1_mid_1 = 1'b0;
			end
		BINARY_223:
			begin
			force_valid_1_2_top_2 = neighbor_force_valid_1[1];
			force_valid_1_2_mid_2 = 1'b0;
			force_valid_1_3_bottom_1 = 1'b0;
			force_valid_1_3_mid_1 = 1'b0;
			force_valid_1_3_top_1 = 1'b0;
			force_valid_2_1_bottom_1 = 1'b0;
			force_valid_2_1_mid_1 = 1'b0;
			end
		BINARY_231:
			begin
			force_valid_1_3_bottom_1 = neighbor_force_valid_1[1];
			force_valid_1_2_mid_2 = 1'b0;
			force_valid_1_2_top_2 = 1'b0;
			force_valid_1_3_mid_1 = 1'b0;
			force_valid_1_3_top_1 = 1'b0;
			force_valid_2_1_bottom_1 = 1'b0;
			force_valid_2_1_mid_1 = 1'b0;
			end
		BINARY_232:
			begin
			force_valid_1_3_mid_1 = neighbor_force_valid_1[1];
			force_valid_1_2_mid_2 = 1'b0;
			force_valid_1_2_top_2 = 1'b0;
			force_valid_1_3_bottom_1 = 1'b0;
			force_valid_1_3_top_1 = 1'b0;
			force_valid_2_1_bottom_1 = 1'b0;
			force_valid_2_1_mid_1 = 1'b0;
			end
		BINARY_233:
			begin
			force_valid_1_3_top_1 = neighbor_force_valid_1[1];
			force_valid_1_2_mid_2 = 1'b0;
			force_valid_1_2_top_2 = 1'b0;
			force_valid_1_3_bottom_1 = 1'b0;
			force_valid_1_3_mid_1 = 1'b0;
			force_valid_2_1_bottom_1 = 1'b0;
			force_valid_2_1_mid_1 = 1'b0;
			end
		BINARY_311:
			begin
			force_valid_2_1_bottom_1 = neighbor_force_valid_1[1];
			force_valid_1_2_mid_2 = 1'b0;
			force_valid_1_2_top_2 = 1'b0;
			force_valid_1_3_bottom_1 = 1'b0;
			force_valid_1_3_mid_1 = 1'b0;
			force_valid_1_3_top_1 = 1'b0;
			force_valid_2_1_mid_1 = 1'b0;
			end
		BINARY_312:
			begin
			force_valid_2_1_mid_1 = neighbor_force_valid_1[1];
			force_valid_1_2_mid_2 = 1'b0;
			force_valid_1_2_top_2 = 1'b0;
			force_valid_1_3_bottom_1 = 1'b0;
			force_valid_1_3_mid_1 = 1'b0;
			force_valid_1_3_top_1 = 1'b0;
			force_valid_2_1_bottom_1 = 1'b0;
			end
		default:
			begin
			force_valid_1_2_mid_2 = 1'b0;
			force_valid_1_2_top_2 = 1'b0;
			force_valid_1_3_bottom_1 = 1'b0;
			force_valid_1_3_mid_1 = 1'b0;
			force_valid_1_3_top_1 = 1'b0;
			force_valid_2_1_bottom_1 = 1'b0;
			force_valid_2_1_mid_1 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_1[2*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:2*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_222:
			begin
			force_valid_1_3_mid_2 = neighbor_force_valid_1[2];
			force_valid_1_3_top_2 = 1'b0;
			force_valid_1_4_bottom_1 = 1'b0;
			force_valid_1_4_mid_1 = 1'b0;
			force_valid_1_4_top_1 = 1'b0;
			force_valid_2_2_bottom_1 = 1'b0;
			force_valid_2_2_mid_1 = 1'b0;
			end
		BINARY_223:
			begin
			force_valid_1_3_top_2 = neighbor_force_valid_1[2];
			force_valid_1_3_mid_2 = 1'b0;
			force_valid_1_4_bottom_1 = 1'b0;
			force_valid_1_4_mid_1 = 1'b0;
			force_valid_1_4_top_1 = 1'b0;
			force_valid_2_2_bottom_1 = 1'b0;
			force_valid_2_2_mid_1 = 1'b0;
			end
		BINARY_231:
			begin
			force_valid_1_4_bottom_1 = neighbor_force_valid_1[2];
			force_valid_1_3_mid_2 = 1'b0;
			force_valid_1_3_top_2 = 1'b0;
			force_valid_1_4_mid_1 = 1'b0;
			force_valid_1_4_top_1 = 1'b0;
			force_valid_2_2_bottom_1 = 1'b0;
			force_valid_2_2_mid_1 = 1'b0;
			end
		BINARY_232:
			begin
			force_valid_1_4_mid_1 = neighbor_force_valid_1[2];
			force_valid_1_3_mid_2 = 1'b0;
			force_valid_1_3_top_2 = 1'b0;
			force_valid_1_4_bottom_1 = 1'b0;
			force_valid_1_4_top_1 = 1'b0;
			force_valid_2_2_bottom_1 = 1'b0;
			force_valid_2_2_mid_1 = 1'b0;
			end
		BINARY_233:
			begin
			force_valid_1_4_top_1 = neighbor_force_valid_1[2];
			force_valid_1_3_mid_2 = 1'b0;
			force_valid_1_3_top_2 = 1'b0;
			force_valid_1_4_bottom_1 = 1'b0;
			force_valid_1_4_mid_1 = 1'b0;
			force_valid_2_2_bottom_1 = 1'b0;
			force_valid_2_2_mid_1 = 1'b0;
			end
		BINARY_311:
			begin
			force_valid_2_2_bottom_1 = neighbor_force_valid_1[2];
			force_valid_1_3_mid_2 = 1'b0;
			force_valid_1_3_top_2 = 1'b0;
			force_valid_1_4_bottom_1 = 1'b0;
			force_valid_1_4_mid_1 = 1'b0;
			force_valid_1_4_top_1 = 1'b0;
			force_valid_2_2_mid_1 = 1'b0;
			end
		BINARY_312:
			begin
			force_valid_2_2_mid_1 = neighbor_force_valid_1[2];
			force_valid_1_3_mid_2 = 1'b0;
			force_valid_1_3_top_2 = 1'b0;
			force_valid_1_4_bottom_1 = 1'b0;
			force_valid_1_4_mid_1 = 1'b0;
			force_valid_1_4_top_1 = 1'b0;
			force_valid_2_2_bottom_1 = 1'b0;
			end
		default:
			begin
			force_valid_1_3_mid_2 = 1'b0;
			force_valid_1_3_top_2 = 1'b0;
			force_valid_1_4_bottom_1 = 1'b0;
			force_valid_1_4_mid_1 = 1'b0;
			force_valid_1_4_top_1 = 1'b0;
			force_valid_2_2_bottom_1 = 1'b0;
			force_valid_2_2_mid_1 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_1[3*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:3*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_222:
			begin
			force_valid_1_4_mid_2 = neighbor_force_valid_1[3];
			force_valid_1_4_top_2 = 1'b0;
			force_valid_1_1_bottom_1 = 1'b0;
			force_valid_1_1_mid_2 = 1'b0;
			force_valid_1_1_top_2 = 1'b0;
			force_valid_2_3_bottom_1 = 1'b0;
			force_valid_2_3_mid_1 = 1'b0;
			end
		BINARY_223:
			begin
			force_valid_1_4_top_2 = neighbor_force_valid_1[3];
			force_valid_1_4_mid_2 = 1'b0;
			force_valid_1_1_bottom_1 = 1'b0;
			force_valid_1_1_mid_2 = 1'b0;
			force_valid_1_1_top_2 = 1'b0;
			force_valid_2_3_bottom_1 = 1'b0;
			force_valid_2_3_mid_1 = 1'b0;
			end
		BINARY_231:
			begin
			force_valid_1_1_bottom_1 = neighbor_force_valid_1[3];
			force_valid_1_4_mid_2 = 1'b0;
			force_valid_1_4_top_2 = 1'b0;
			force_valid_1_1_mid_2 = 1'b0;
			force_valid_1_1_top_2 = 1'b0;
			force_valid_2_3_bottom_1 = 1'b0;
			force_valid_2_3_mid_1 = 1'b0;
			end
		BINARY_232:
			begin
			force_valid_1_1_mid_2 = neighbor_force_valid_1[3];
			force_valid_1_4_mid_2 = 1'b0;
			force_valid_1_4_top_2 = 1'b0;
			force_valid_1_1_bottom_1 = 1'b0;
			force_valid_1_1_top_2 = 1'b0;
			force_valid_2_3_bottom_1 = 1'b0;
			force_valid_2_3_mid_1 = 1'b0;
			end
		BINARY_233:
			begin
			force_valid_1_1_top_2 = neighbor_force_valid_1[3];
			force_valid_1_4_mid_2 = 1'b0;
			force_valid_1_4_top_2 = 1'b0;
			force_valid_1_1_bottom_1 = 1'b0;
			force_valid_1_1_mid_2 = 1'b0;
			force_valid_2_3_bottom_1 = 1'b0;
			force_valid_2_3_mid_1 = 1'b0;
			end
		BINARY_311:
			begin
			force_valid_2_3_bottom_1 = neighbor_force_valid_1[3];
			force_valid_1_4_mid_2 = 1'b0;
			force_valid_1_4_top_2 = 1'b0;
			force_valid_1_1_bottom_1 = 1'b0;
			force_valid_1_1_mid_2 = 1'b0;
			force_valid_1_1_top_2 = 1'b0;
			force_valid_2_3_mid_1 = 1'b0;
			end
		BINARY_312:
			begin
			force_valid_2_3_mid_1 = neighbor_force_valid_1[3];
			force_valid_1_4_mid_2 = 1'b0;
			force_valid_1_4_top_2 = 1'b0;
			force_valid_1_1_bottom_1 = 1'b0;
			force_valid_1_1_mid_2 = 1'b0;
			force_valid_1_1_top_2 = 1'b0;
			force_valid_2_3_bottom_1 = 1'b0;
			end
		default:
			begin
			force_valid_1_4_mid_2 = 1'b0;
			force_valid_1_4_top_2 = 1'b0;
			force_valid_1_1_bottom_1 = 1'b0;
			force_valid_1_1_mid_2 = 1'b0;
			force_valid_1_1_top_2 = 1'b0;
			force_valid_2_3_bottom_1 = 1'b0;
			force_valid_2_3_mid_1 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_1[4*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:4*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_222:
			begin
			force_valid_2_1_mid_2 = neighbor_force_valid_1[4];
			force_valid_2_1_top_1 = 1'b0;
			force_valid_2_2_bottom_2 = 1'b0;
			force_valid_2_2_mid_2 = 1'b0;
			force_valid_2_2_top_1 = 1'b0;
			force_valid_3_4_bottom_1 = 1'b0;
			force_valid_3_4_mid_1 = 1'b0;
			end
		BINARY_223:
			begin
			force_valid_2_1_top_1 = neighbor_force_valid_1[4];
			force_valid_2_1_mid_2 = 1'b0;
			force_valid_2_2_bottom_2 = 1'b0;
			force_valid_2_2_mid_2 = 1'b0;
			force_valid_2_2_top_1 = 1'b0;
			force_valid_3_4_bottom_1 = 1'b0;
			force_valid_3_4_mid_1 = 1'b0;
			end
		BINARY_231:
			begin
			force_valid_2_2_bottom_2 = neighbor_force_valid_1[4];
			force_valid_2_1_mid_2 = 1'b0;
			force_valid_2_1_top_1 = 1'b0;
			force_valid_2_2_mid_2 = 1'b0;
			force_valid_2_2_top_1 = 1'b0;
			force_valid_3_4_bottom_1 = 1'b0;
			force_valid_3_4_mid_1 = 1'b0;
			end
		BINARY_232:
			begin
			force_valid_2_2_mid_2 = neighbor_force_valid_1[4];
			force_valid_2_1_mid_2 = 1'b0;
			force_valid_2_1_top_1 = 1'b0;
			force_valid_2_2_bottom_2 = 1'b0;
			force_valid_2_2_top_1 = 1'b0;
			force_valid_3_4_bottom_1 = 1'b0;
			force_valid_3_4_mid_1 = 1'b0;
			end
		BINARY_233:
			begin
			force_valid_2_2_top_1 = neighbor_force_valid_1[4];
			force_valid_2_1_mid_2 = 1'b0;
			force_valid_2_1_top_1 = 1'b0;
			force_valid_2_2_bottom_2 = 1'b0;
			force_valid_2_2_mid_2 = 1'b0;
			force_valid_3_4_bottom_1 = 1'b0;
			force_valid_3_4_mid_1 = 1'b0;
			end
		BINARY_311:
			begin
			force_valid_3_4_bottom_1 = neighbor_force_valid_1[4];
			force_valid_2_1_mid_2 = 1'b0;
			force_valid_2_1_top_1 = 1'b0;
			force_valid_2_2_bottom_2 = 1'b0;
			force_valid_2_2_mid_2 = 1'b0;
			force_valid_2_2_top_1 = 1'b0;
			force_valid_3_4_mid_1 = 1'b0;
			end
		BINARY_312:
			begin
			force_valid_3_4_mid_1 = neighbor_force_valid_1[4];
			force_valid_2_1_mid_2 = 1'b0;
			force_valid_2_1_top_1 = 1'b0;
			force_valid_2_2_bottom_2 = 1'b0;
			force_valid_2_2_mid_2 = 1'b0;
			force_valid_2_2_top_1 = 1'b0;
			force_valid_3_4_bottom_1 = 1'b0;
			end
		default:
			begin
			force_valid_2_1_mid_2 = 1'b0;
			force_valid_2_1_top_1 = 1'b0;
			force_valid_2_2_bottom_2 = 1'b0;
			force_valid_2_2_mid_2 = 1'b0;
			force_valid_2_2_top_1 = 1'b0;
			force_valid_3_4_bottom_1 = 1'b0;
			force_valid_3_4_mid_1 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_1[5*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:5*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_222:
			begin
			force_valid_2_2_mid_3 = neighbor_force_valid_1[5];
			force_valid_2_2_top_2 = 1'b0;
			force_valid_2_3_bottom_2 = 1'b0;
			force_valid_2_3_mid_2 = 1'b0;
			force_valid_2_3_top_1 = 1'b0;
			force_valid_3_1_bottom_1 = 1'b0;
			force_valid_3_1_mid_1 = 1'b0;
			end
		BINARY_223:
			begin
			force_valid_2_2_top_2 = neighbor_force_valid_1[5];
			force_valid_2_2_mid_3 = 1'b0;
			force_valid_2_3_bottom_2 = 1'b0;
			force_valid_2_3_mid_2 = 1'b0;
			force_valid_2_3_top_1 = 1'b0;
			force_valid_3_1_bottom_1 = 1'b0;
			force_valid_3_1_mid_1 = 1'b0;
			end
		BINARY_231:
			begin
			force_valid_2_3_bottom_2 = neighbor_force_valid_1[5];
			force_valid_2_2_mid_3 = 1'b0;
			force_valid_2_2_top_2 = 1'b0;
			force_valid_2_3_mid_2 = 1'b0;
			force_valid_2_3_top_1 = 1'b0;
			force_valid_3_1_bottom_1 = 1'b0;
			force_valid_3_1_mid_1 = 1'b0;
			end
		BINARY_232:
			begin
			force_valid_2_3_mid_2 = neighbor_force_valid_1[5];
			force_valid_2_2_mid_3 = 1'b0;
			force_valid_2_2_top_2 = 1'b0;
			force_valid_2_3_bottom_2 = 1'b0;
			force_valid_2_3_top_1 = 1'b0;
			force_valid_3_1_bottom_1 = 1'b0;
			force_valid_3_1_mid_1 = 1'b0;
			end
		BINARY_233:
			begin
			force_valid_2_3_top_1 = neighbor_force_valid_1[5];
			force_valid_2_2_mid_3 = 1'b0;
			force_valid_2_2_top_2 = 1'b0;
			force_valid_2_3_bottom_2 = 1'b0;
			force_valid_2_3_mid_2 = 1'b0;
			force_valid_3_1_bottom_1 = 1'b0;
			force_valid_3_1_mid_1 = 1'b0;
			end
		BINARY_311:
			begin
			force_valid_3_1_bottom_1 = neighbor_force_valid_1[5];
			force_valid_2_2_mid_3 = 1'b0;
			force_valid_2_2_top_2 = 1'b0;
			force_valid_2_3_bottom_2 = 1'b0;
			force_valid_2_3_mid_2 = 1'b0;
			force_valid_2_3_top_1 = 1'b0;
			force_valid_3_1_mid_1 = 1'b0;
			end
		BINARY_312:
			begin
			force_valid_3_1_mid_1 = neighbor_force_valid_1[5];
			force_valid_2_2_mid_3 = 1'b0;
			force_valid_2_2_top_2 = 1'b0;
			force_valid_2_3_bottom_2 = 1'b0;
			force_valid_2_3_mid_2 = 1'b0;
			force_valid_2_3_top_1 = 1'b0;
			force_valid_3_1_bottom_1 = 1'b0;
			end
		default:
			begin
			force_valid_2_2_mid_3 = 1'b0;
			force_valid_2_2_top_2 = 1'b0;
			force_valid_2_3_bottom_2 = 1'b0;
			force_valid_2_3_mid_2 = 1'b0;
			force_valid_2_3_top_1 = 1'b0;
			force_valid_3_1_bottom_1 = 1'b0;
			force_valid_3_1_mid_1 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_1[6*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:6*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_222:
			begin
			force_valid_2_3_mid_3 = neighbor_force_valid_1[6];
			force_valid_2_3_top_2 = 1'b0;
			force_valid_2_4_bottom_2 = 1'b0;
			force_valid_2_4_mid_2 = 1'b0;
			force_valid_2_4_top_1 = 1'b0;
			force_valid_3_2_bottom_1 = 1'b0;
			force_valid_3_2_mid_1 = 1'b0;
			end
		BINARY_223:
			begin
			force_valid_2_3_top_2 = neighbor_force_valid_1[6];
			force_valid_2_3_mid_3 = 1'b0;
			force_valid_2_4_bottom_2 = 1'b0;
			force_valid_2_4_mid_2 = 1'b0;
			force_valid_2_4_top_1 = 1'b0;
			force_valid_3_2_bottom_1 = 1'b0;
			force_valid_3_2_mid_1 = 1'b0;
			end
		BINARY_231:
			begin
			force_valid_2_4_bottom_2 = neighbor_force_valid_1[6];
			force_valid_2_3_mid_3 = 1'b0;
			force_valid_2_3_top_2 = 1'b0;
			force_valid_2_4_mid_2 = 1'b0;
			force_valid_2_4_top_1 = 1'b0;
			force_valid_3_2_bottom_1 = 1'b0;
			force_valid_3_2_mid_1 = 1'b0;
			end
		BINARY_232:
			begin
			force_valid_2_4_mid_2 = neighbor_force_valid_1[6];
			force_valid_2_3_mid_3 = 1'b0;
			force_valid_2_3_top_2 = 1'b0;
			force_valid_2_4_bottom_2 = 1'b0;
			force_valid_2_4_top_1 = 1'b0;
			force_valid_3_2_bottom_1 = 1'b0;
			force_valid_3_2_mid_1 = 1'b0;
			end
		BINARY_233:
			begin
			force_valid_2_4_top_1 = neighbor_force_valid_1[6];
			force_valid_2_3_mid_3 = 1'b0;
			force_valid_2_3_top_2 = 1'b0;
			force_valid_2_4_bottom_2 = 1'b0;
			force_valid_2_4_mid_2 = 1'b0;
			force_valid_3_2_bottom_1 = 1'b0;
			force_valid_3_2_mid_1 = 1'b0;
			end
		BINARY_311:
			begin
			force_valid_3_2_bottom_1 = neighbor_force_valid_1[6];
			force_valid_2_3_mid_3 = 1'b0;
			force_valid_2_3_top_2 = 1'b0;
			force_valid_2_4_bottom_2 = 1'b0;
			force_valid_2_4_mid_2 = 1'b0;
			force_valid_2_4_top_1 = 1'b0;
			force_valid_3_2_mid_1 = 1'b0;
			end
		BINARY_312:
			begin
			force_valid_3_2_mid_1 = neighbor_force_valid_1[6];
			force_valid_2_3_mid_3 = 1'b0;
			force_valid_2_3_top_2 = 1'b0;
			force_valid_2_4_bottom_2 = 1'b0;
			force_valid_2_4_mid_2 = 1'b0;
			force_valid_2_4_top_1 = 1'b0;
			force_valid_3_2_bottom_1 = 1'b0;
			end
		default:
			begin
			force_valid_2_3_mid_3 = 1'b0;
			force_valid_2_3_top_2 = 1'b0;
			force_valid_2_4_bottom_2 = 1'b0;
			force_valid_2_4_mid_2 = 1'b0;
			force_valid_2_4_top_1 = 1'b0;
			force_valid_3_2_bottom_1 = 1'b0;
			force_valid_3_2_mid_1 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_1[7*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:7*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_222:
			begin
			force_valid_2_4_mid_3 = neighbor_force_valid_1[7];
			force_valid_2_4_top_2 = 1'b0;
			force_valid_2_1_bottom_2 = 1'b0;
			force_valid_2_1_mid_3 = 1'b0;
			force_valid_2_1_top_2 = 1'b0;
			force_valid_3_3_bottom_1 = 1'b0;
			force_valid_3_3_mid_1 = 1'b0;
			end
		BINARY_223:
			begin
			force_valid_2_4_top_2 = neighbor_force_valid_1[7];
			force_valid_2_4_mid_3 = 1'b0;
			force_valid_2_1_bottom_2 = 1'b0;
			force_valid_2_1_mid_3 = 1'b0;
			force_valid_2_1_top_2 = 1'b0;
			force_valid_3_3_bottom_1 = 1'b0;
			force_valid_3_3_mid_1 = 1'b0;
			end
		BINARY_231:
			begin
			force_valid_2_1_bottom_2 = neighbor_force_valid_1[7];
			force_valid_2_4_mid_3 = 1'b0;
			force_valid_2_4_top_2 = 1'b0;
			force_valid_2_1_mid_3 = 1'b0;
			force_valid_2_1_top_2 = 1'b0;
			force_valid_3_3_bottom_1 = 1'b0;
			force_valid_3_3_mid_1 = 1'b0;
			end
		BINARY_232:
			begin
			force_valid_2_1_mid_3 = neighbor_force_valid_1[7];
			force_valid_2_4_mid_3 = 1'b0;
			force_valid_2_4_top_2 = 1'b0;
			force_valid_2_1_bottom_2 = 1'b0;
			force_valid_2_1_top_2 = 1'b0;
			force_valid_3_3_bottom_1 = 1'b0;
			force_valid_3_3_mid_1 = 1'b0;
			end
		BINARY_233:
			begin
			force_valid_2_1_top_2 = neighbor_force_valid_1[7];
			force_valid_2_4_mid_3 = 1'b0;
			force_valid_2_4_top_2 = 1'b0;
			force_valid_2_1_bottom_2 = 1'b0;
			force_valid_2_1_mid_3 = 1'b0;
			force_valid_3_3_bottom_1 = 1'b0;
			force_valid_3_3_mid_1 = 1'b0;
			end
		BINARY_311:
			begin
			force_valid_3_3_bottom_1 = neighbor_force_valid_1[7];
			force_valid_2_4_mid_3 = 1'b0;
			force_valid_2_4_top_2 = 1'b0;
			force_valid_2_1_bottom_2 = 1'b0;
			force_valid_2_1_mid_3 = 1'b0;
			force_valid_2_1_top_2 = 1'b0;
			force_valid_3_3_mid_1 = 1'b0;
			end
		BINARY_312:
			begin
			force_valid_3_3_mid_1 = neighbor_force_valid_1[7];
			force_valid_2_4_mid_3 = 1'b0;
			force_valid_2_4_top_2 = 1'b0;
			force_valid_2_1_bottom_2 = 1'b0;
			force_valid_2_1_mid_3 = 1'b0;
			force_valid_2_1_top_2 = 1'b0;
			force_valid_3_3_bottom_1 = 1'b0;
			end
		default:
			begin
			force_valid_2_4_mid_3 = 1'b0;
			force_valid_2_4_top_2 = 1'b0;
			force_valid_2_1_bottom_2 = 1'b0;
			force_valid_2_1_mid_3 = 1'b0;
			force_valid_2_1_top_2 = 1'b0;
			force_valid_3_3_bottom_1 = 1'b0;
			force_valid_3_3_mid_1 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_1[8*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:8*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_222:
			begin
			force_valid_3_1_mid_2 = neighbor_force_valid_1[8];
			force_valid_3_1_top_1 = 1'b0;
			force_valid_3_2_bottom_2 = 1'b0;
			force_valid_3_2_mid_2 = 1'b0;
			force_valid_3_2_top_1 = 1'b0;
			force_valid_4_4_bottom_1 = 1'b0;
			force_valid_4_4_mid_1 = 1'b0;
			end
		BINARY_223:
			begin
			force_valid_3_1_top_1 = neighbor_force_valid_1[8];
			force_valid_3_1_mid_2 = 1'b0;
			force_valid_3_2_bottom_2 = 1'b0;
			force_valid_3_2_mid_2 = 1'b0;
			force_valid_3_2_top_1 = 1'b0;
			force_valid_4_4_bottom_1 = 1'b0;
			force_valid_4_4_mid_1 = 1'b0;
			end
		BINARY_231:
			begin
			force_valid_3_2_bottom_2 = neighbor_force_valid_1[8];
			force_valid_3_1_mid_2 = 1'b0;
			force_valid_3_1_top_1 = 1'b0;
			force_valid_3_2_mid_2 = 1'b0;
			force_valid_3_2_top_1 = 1'b0;
			force_valid_4_4_bottom_1 = 1'b0;
			force_valid_4_4_mid_1 = 1'b0;
			end
		BINARY_232:
			begin
			force_valid_3_2_mid_2 = neighbor_force_valid_1[8];
			force_valid_3_1_mid_2 = 1'b0;
			force_valid_3_1_top_1 = 1'b0;
			force_valid_3_2_bottom_2 = 1'b0;
			force_valid_3_2_top_1 = 1'b0;
			force_valid_4_4_bottom_1 = 1'b0;
			force_valid_4_4_mid_1 = 1'b0;
			end
		BINARY_233:
			begin
			force_valid_3_2_top_1 = neighbor_force_valid_1[8];
			force_valid_3_1_mid_2 = 1'b0;
			force_valid_3_1_top_1 = 1'b0;
			force_valid_3_2_bottom_2 = 1'b0;
			force_valid_3_2_mid_2 = 1'b0;
			force_valid_4_4_bottom_1 = 1'b0;
			force_valid_4_4_mid_1 = 1'b0;
			end
		BINARY_311:
			begin
			force_valid_4_4_bottom_1 = neighbor_force_valid_1[8];
			force_valid_3_1_mid_2 = 1'b0;
			force_valid_3_1_top_1 = 1'b0;
			force_valid_3_2_bottom_2 = 1'b0;
			force_valid_3_2_mid_2 = 1'b0;
			force_valid_3_2_top_1 = 1'b0;
			force_valid_4_4_mid_1 = 1'b0;
			end
		BINARY_312:
			begin
			force_valid_4_4_mid_1 = neighbor_force_valid_1[8];
			force_valid_3_1_mid_2 = 1'b0;
			force_valid_3_1_top_1 = 1'b0;
			force_valid_3_2_bottom_2 = 1'b0;
			force_valid_3_2_mid_2 = 1'b0;
			force_valid_3_2_top_1 = 1'b0;
			force_valid_4_4_bottom_1 = 1'b0;
			end
		default:
			begin
			force_valid_3_1_mid_2 = 1'b0;
			force_valid_3_1_top_1 = 1'b0;
			force_valid_3_2_bottom_2 = 1'b0;
			force_valid_3_2_mid_2 = 1'b0;
			force_valid_3_2_top_1 = 1'b0;
			force_valid_4_4_bottom_1 = 1'b0;
			force_valid_4_4_mid_1 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_1[9*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:9*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_222:
			begin
			force_valid_3_2_mid_3 = neighbor_force_valid_1[9];
			force_valid_3_2_top_2 = 1'b0;
			force_valid_3_3_bottom_2 = 1'b0;
			force_valid_3_3_mid_2 = 1'b0;
			force_valid_3_3_top_1 = 1'b0;
			force_valid_4_1_bottom_1 = 1'b0;
			force_valid_4_1_mid_1 = 1'b0;
			end
		BINARY_223:
			begin
			force_valid_3_2_top_2 = neighbor_force_valid_1[9];
			force_valid_3_2_mid_3 = 1'b0;
			force_valid_3_3_bottom_2 = 1'b0;
			force_valid_3_3_mid_2 = 1'b0;
			force_valid_3_3_top_1 = 1'b0;
			force_valid_4_1_bottom_1 = 1'b0;
			force_valid_4_1_mid_1 = 1'b0;
			end
		BINARY_231:
			begin
			force_valid_3_3_bottom_2 = neighbor_force_valid_1[9];
			force_valid_3_2_mid_3 = 1'b0;
			force_valid_3_2_top_2 = 1'b0;
			force_valid_3_3_mid_2 = 1'b0;
			force_valid_3_3_top_1 = 1'b0;
			force_valid_4_1_bottom_1 = 1'b0;
			force_valid_4_1_mid_1 = 1'b0;
			end
		BINARY_232:
			begin
			force_valid_3_3_mid_2 = neighbor_force_valid_1[9];
			force_valid_3_2_mid_3 = 1'b0;
			force_valid_3_2_top_2 = 1'b0;
			force_valid_3_3_bottom_2 = 1'b0;
			force_valid_3_3_top_1 = 1'b0;
			force_valid_4_1_bottom_1 = 1'b0;
			force_valid_4_1_mid_1 = 1'b0;
			end
		BINARY_233:
			begin
			force_valid_3_3_top_1 = neighbor_force_valid_1[9];
			force_valid_3_2_mid_3 = 1'b0;
			force_valid_3_2_top_2 = 1'b0;
			force_valid_3_3_bottom_2 = 1'b0;
			force_valid_3_3_mid_2 = 1'b0;
			force_valid_4_1_bottom_1 = 1'b0;
			force_valid_4_1_mid_1 = 1'b0;
			end
		BINARY_311:
			begin
			force_valid_4_1_bottom_1 = neighbor_force_valid_1[9];
			force_valid_3_2_mid_3 = 1'b0;
			force_valid_3_2_top_2 = 1'b0;
			force_valid_3_3_bottom_2 = 1'b0;
			force_valid_3_3_mid_2 = 1'b0;
			force_valid_3_3_top_1 = 1'b0;
			force_valid_4_1_mid_1 = 1'b0;
			end
		BINARY_312:
			begin
			force_valid_4_1_mid_1 = neighbor_force_valid_1[9];
			force_valid_3_2_mid_3 = 1'b0;
			force_valid_3_2_top_2 = 1'b0;
			force_valid_3_3_bottom_2 = 1'b0;
			force_valid_3_3_mid_2 = 1'b0;
			force_valid_3_3_top_1 = 1'b0;
			force_valid_4_1_bottom_1 = 1'b0;
			end
		default:
			begin
			force_valid_3_2_mid_3 = 1'b0;
			force_valid_3_2_top_2 = 1'b0;
			force_valid_3_3_bottom_2 = 1'b0;
			force_valid_3_3_mid_2 = 1'b0;
			force_valid_3_3_top_1 = 1'b0;
			force_valid_4_1_bottom_1 = 1'b0;
			force_valid_4_1_mid_1 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_1[10*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:10*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_222:
			begin
			force_valid_3_3_mid_3 = neighbor_force_valid_1[10];
			force_valid_3_3_top_2 = 1'b0;
			force_valid_3_4_bottom_2 = 1'b0;
			force_valid_3_4_mid_2 = 1'b0;
			force_valid_3_4_top_1 = 1'b0;
			force_valid_4_2_bottom_1 = 1'b0;
			force_valid_4_2_mid_1 = 1'b0;
			end
		BINARY_223:
			begin
			force_valid_3_3_top_2 = neighbor_force_valid_1[10];
			force_valid_3_3_mid_3 = 1'b0;
			force_valid_3_4_bottom_2 = 1'b0;
			force_valid_3_4_mid_2 = 1'b0;
			force_valid_3_4_top_1 = 1'b0;
			force_valid_4_2_bottom_1 = 1'b0;
			force_valid_4_2_mid_1 = 1'b0;
			end
		BINARY_231:
			begin
			force_valid_3_4_bottom_2 = neighbor_force_valid_1[10];
			force_valid_3_3_mid_3 = 1'b0;
			force_valid_3_3_top_2 = 1'b0;
			force_valid_3_4_mid_2 = 1'b0;
			force_valid_3_4_top_1 = 1'b0;
			force_valid_4_2_bottom_1 = 1'b0;
			force_valid_4_2_mid_1 = 1'b0;
			end
		BINARY_232:
			begin
			force_valid_3_4_mid_2 = neighbor_force_valid_1[10];
			force_valid_3_3_mid_3 = 1'b0;
			force_valid_3_3_top_2 = 1'b0;
			force_valid_3_4_bottom_2 = 1'b0;
			force_valid_3_4_top_1 = 1'b0;
			force_valid_4_2_bottom_1 = 1'b0;
			force_valid_4_2_mid_1 = 1'b0;
			end
		BINARY_233:
			begin
			force_valid_3_4_top_1 = neighbor_force_valid_1[10];
			force_valid_3_3_mid_3 = 1'b0;
			force_valid_3_3_top_2 = 1'b0;
			force_valid_3_4_bottom_2 = 1'b0;
			force_valid_3_4_mid_2 = 1'b0;
			force_valid_4_2_bottom_1 = 1'b0;
			force_valid_4_2_mid_1 = 1'b0;
			end
		BINARY_311:
			begin
			force_valid_4_2_bottom_1 = neighbor_force_valid_1[10];
			force_valid_3_3_mid_3 = 1'b0;
			force_valid_3_3_top_2 = 1'b0;
			force_valid_3_4_bottom_2 = 1'b0;
			force_valid_3_4_mid_2 = 1'b0;
			force_valid_3_4_top_1 = 1'b0;
			force_valid_4_2_mid_1 = 1'b0;
			end
		BINARY_312:
			begin
			force_valid_4_2_mid_1 = neighbor_force_valid_1[10];
			force_valid_3_3_mid_3 = 1'b0;
			force_valid_3_3_top_2 = 1'b0;
			force_valid_3_4_bottom_2 = 1'b0;
			force_valid_3_4_mid_2 = 1'b0;
			force_valid_3_4_top_1 = 1'b0;
			force_valid_4_2_bottom_1 = 1'b0;
			end
		default:
			begin
			force_valid_3_3_mid_3 = 1'b0;
			force_valid_3_3_top_2 = 1'b0;
			force_valid_3_4_bottom_2 = 1'b0;
			force_valid_3_4_mid_2 = 1'b0;
			force_valid_3_4_top_1 = 1'b0;
			force_valid_4_2_bottom_1 = 1'b0;
			force_valid_4_2_mid_1 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_1[11*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:11*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_222:
			begin
			force_valid_3_4_mid_3 = neighbor_force_valid_1[11];
			force_valid_3_4_top_2 = 1'b0;
			force_valid_3_1_bottom_2 = 1'b0;
			force_valid_3_1_mid_3 = 1'b0;
			force_valid_3_1_top_2 = 1'b0;
			force_valid_4_3_bottom_1 = 1'b0;
			force_valid_4_3_mid_1 = 1'b0;
			end
		BINARY_223:
			begin
			force_valid_3_4_top_2 = neighbor_force_valid_1[11];
			force_valid_3_4_mid_3 = 1'b0;
			force_valid_3_1_bottom_2 = 1'b0;
			force_valid_3_1_mid_3 = 1'b0;
			force_valid_3_1_top_2 = 1'b0;
			force_valid_4_3_bottom_1 = 1'b0;
			force_valid_4_3_mid_1 = 1'b0;
			end
		BINARY_231:
			begin
			force_valid_3_1_bottom_2 = neighbor_force_valid_1[11];
			force_valid_3_4_mid_3 = 1'b0;
			force_valid_3_4_top_2 = 1'b0;
			force_valid_3_1_mid_3 = 1'b0;
			force_valid_3_1_top_2 = 1'b0;
			force_valid_4_3_bottom_1 = 1'b0;
			force_valid_4_3_mid_1 = 1'b0;
			end
		BINARY_232:
			begin
			force_valid_3_1_mid_3 = neighbor_force_valid_1[11];
			force_valid_3_4_mid_3 = 1'b0;
			force_valid_3_4_top_2 = 1'b0;
			force_valid_3_1_bottom_2 = 1'b0;
			force_valid_3_1_top_2 = 1'b0;
			force_valid_4_3_bottom_1 = 1'b0;
			force_valid_4_3_mid_1 = 1'b0;
			end
		BINARY_233:
			begin
			force_valid_3_1_top_2 = neighbor_force_valid_1[11];
			force_valid_3_4_mid_3 = 1'b0;
			force_valid_3_4_top_2 = 1'b0;
			force_valid_3_1_bottom_2 = 1'b0;
			force_valid_3_1_mid_3 = 1'b0;
			force_valid_4_3_bottom_1 = 1'b0;
			force_valid_4_3_mid_1 = 1'b0;
			end
		BINARY_311:
			begin
			force_valid_4_3_bottom_1 = neighbor_force_valid_1[11];
			force_valid_3_4_mid_3 = 1'b0;
			force_valid_3_4_top_2 = 1'b0;
			force_valid_3_1_bottom_2 = 1'b0;
			force_valid_3_1_mid_3 = 1'b0;
			force_valid_3_1_top_2 = 1'b0;
			force_valid_4_3_mid_1 = 1'b0;
			end
		BINARY_312:
			begin
			force_valid_4_3_mid_1 = neighbor_force_valid_1[11];
			force_valid_3_4_mid_3 = 1'b0;
			force_valid_3_4_top_2 = 1'b0;
			force_valid_3_1_bottom_2 = 1'b0;
			force_valid_3_1_mid_3 = 1'b0;
			force_valid_3_1_top_2 = 1'b0;
			force_valid_4_3_bottom_1 = 1'b0;
			end
		default:
			begin
			force_valid_3_4_mid_3 = 1'b0;
			force_valid_3_4_top_2 = 1'b0;
			force_valid_3_1_bottom_2 = 1'b0;
			force_valid_3_1_mid_3 = 1'b0;
			force_valid_3_1_top_2 = 1'b0;
			force_valid_4_3_bottom_1 = 1'b0;
			force_valid_4_3_mid_1 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_1[12*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:12*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_222:
			begin
			force_valid_4_1_mid_2 = neighbor_force_valid_1[12];
			force_valid_4_1_top_1 = 1'b0;
			force_valid_4_2_bottom_2 = 1'b0;
			force_valid_4_2_mid_2 = 1'b0;
			force_valid_4_2_top_1 = 1'b0;
			force_valid_1_4_bottom_2 = 1'b0;
			force_valid_1_4_mid_3 = 1'b0;
			end
		BINARY_223:
			begin
			force_valid_4_1_top_1 = neighbor_force_valid_1[12];
			force_valid_4_1_mid_2 = 1'b0;
			force_valid_4_2_bottom_2 = 1'b0;
			force_valid_4_2_mid_2 = 1'b0;
			force_valid_4_2_top_1 = 1'b0;
			force_valid_1_4_bottom_2 = 1'b0;
			force_valid_1_4_mid_3 = 1'b0;
			end
		BINARY_231:
			begin
			force_valid_4_2_bottom_2 = neighbor_force_valid_1[12];
			force_valid_4_1_mid_2 = 1'b0;
			force_valid_4_1_top_1 = 1'b0;
			force_valid_4_2_mid_2 = 1'b0;
			force_valid_4_2_top_1 = 1'b0;
			force_valid_1_4_bottom_2 = 1'b0;
			force_valid_1_4_mid_3 = 1'b0;
			end
		BINARY_232:
			begin
			force_valid_4_2_mid_2 = neighbor_force_valid_1[12];
			force_valid_4_1_mid_2 = 1'b0;
			force_valid_4_1_top_1 = 1'b0;
			force_valid_4_2_bottom_2 = 1'b0;
			force_valid_4_2_top_1 = 1'b0;
			force_valid_1_4_bottom_2 = 1'b0;
			force_valid_1_4_mid_3 = 1'b0;
			end
		BINARY_233:
			begin
			force_valid_4_2_top_1 = neighbor_force_valid_1[12];
			force_valid_4_1_mid_2 = 1'b0;
			force_valid_4_1_top_1 = 1'b0;
			force_valid_4_2_bottom_2 = 1'b0;
			force_valid_4_2_mid_2 = 1'b0;
			force_valid_1_4_bottom_2 = 1'b0;
			force_valid_1_4_mid_3 = 1'b0;
			end
		BINARY_311:
			begin
			force_valid_1_4_bottom_2 = neighbor_force_valid_1[12];
			force_valid_4_1_mid_2 = 1'b0;
			force_valid_4_1_top_1 = 1'b0;
			force_valid_4_2_bottom_2 = 1'b0;
			force_valid_4_2_mid_2 = 1'b0;
			force_valid_4_2_top_1 = 1'b0;
			force_valid_1_4_mid_3 = 1'b0;
			end
		BINARY_312:
			begin
			force_valid_1_4_mid_3 = neighbor_force_valid_1[12];
			force_valid_4_1_mid_2 = 1'b0;
			force_valid_4_1_top_1 = 1'b0;
			force_valid_4_2_bottom_2 = 1'b0;
			force_valid_4_2_mid_2 = 1'b0;
			force_valid_4_2_top_1 = 1'b0;
			force_valid_1_4_bottom_2 = 1'b0;
			end
		default:
			begin
			force_valid_4_1_mid_2 = 1'b0;
			force_valid_4_1_top_1 = 1'b0;
			force_valid_4_2_bottom_2 = 1'b0;
			force_valid_4_2_mid_2 = 1'b0;
			force_valid_4_2_top_1 = 1'b0;
			force_valid_1_4_bottom_2 = 1'b0;
			force_valid_1_4_mid_3 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_1[13*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:13*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_222:
			begin
			force_valid_4_2_mid_3 = neighbor_force_valid_1[13];
			force_valid_4_2_top_2 = 1'b0;
			force_valid_4_3_bottom_2 = 1'b0;
			force_valid_4_3_mid_2 = 1'b0;
			force_valid_4_3_top_1 = 1'b0;
			force_valid_1_1_bottom_2 = 1'b0;
			force_valid_1_1_mid_3 = 1'b0;
			end
		BINARY_223:
			begin
			force_valid_4_2_top_2 = neighbor_force_valid_1[13];
			force_valid_4_2_mid_3 = 1'b0;
			force_valid_4_3_bottom_2 = 1'b0;
			force_valid_4_3_mid_2 = 1'b0;
			force_valid_4_3_top_1 = 1'b0;
			force_valid_1_1_bottom_2 = 1'b0;
			force_valid_1_1_mid_3 = 1'b0;
			end
		BINARY_231:
			begin
			force_valid_4_3_bottom_2 = neighbor_force_valid_1[13];
			force_valid_4_2_mid_3 = 1'b0;
			force_valid_4_2_top_2 = 1'b0;
			force_valid_4_3_mid_2 = 1'b0;
			force_valid_4_3_top_1 = 1'b0;
			force_valid_1_1_bottom_2 = 1'b0;
			force_valid_1_1_mid_3 = 1'b0;
			end
		BINARY_232:
			begin
			force_valid_4_3_mid_2 = neighbor_force_valid_1[13];
			force_valid_4_2_mid_3 = 1'b0;
			force_valid_4_2_top_2 = 1'b0;
			force_valid_4_3_bottom_2 = 1'b0;
			force_valid_4_3_top_1 = 1'b0;
			force_valid_1_1_bottom_2 = 1'b0;
			force_valid_1_1_mid_3 = 1'b0;
			end
		BINARY_233:
			begin
			force_valid_4_3_top_1 = neighbor_force_valid_1[13];
			force_valid_4_2_mid_3 = 1'b0;
			force_valid_4_2_top_2 = 1'b0;
			force_valid_4_3_bottom_2 = 1'b0;
			force_valid_4_3_mid_2 = 1'b0;
			force_valid_1_1_bottom_2 = 1'b0;
			force_valid_1_1_mid_3 = 1'b0;
			end
		BINARY_311:
			begin
			force_valid_1_1_bottom_2 = neighbor_force_valid_1[13];
			force_valid_4_2_mid_3 = 1'b0;
			force_valid_4_2_top_2 = 1'b0;
			force_valid_4_3_bottom_2 = 1'b0;
			force_valid_4_3_mid_2 = 1'b0;
			force_valid_4_3_top_1 = 1'b0;
			force_valid_1_1_mid_3 = 1'b0;
			end
		BINARY_312:
			begin
			force_valid_1_1_mid_3 = neighbor_force_valid_1[13];
			force_valid_4_2_mid_3 = 1'b0;
			force_valid_4_2_top_2 = 1'b0;
			force_valid_4_3_bottom_2 = 1'b0;
			force_valid_4_3_mid_2 = 1'b0;
			force_valid_4_3_top_1 = 1'b0;
			force_valid_1_1_bottom_2 = 1'b0;
			end
		default:
			begin
			force_valid_4_2_mid_3 = 1'b0;
			force_valid_4_2_top_2 = 1'b0;
			force_valid_4_3_bottom_2 = 1'b0;
			force_valid_4_3_mid_2 = 1'b0;
			force_valid_4_3_top_1 = 1'b0;
			force_valid_1_1_bottom_2 = 1'b0;
			force_valid_1_1_mid_3 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_1[14*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:14*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_222:
			begin
			force_valid_4_3_mid_3 = neighbor_force_valid_1[14];
			force_valid_4_3_top_2 = 1'b0;
			force_valid_4_4_bottom_2 = 1'b0;
			force_valid_4_4_mid_2 = 1'b0;
			force_valid_4_4_top_1 = 1'b0;
			force_valid_1_2_bottom_2 = 1'b0;
			force_valid_1_2_mid_3 = 1'b0;
			end
		BINARY_223:
			begin
			force_valid_4_3_top_2 = neighbor_force_valid_1[14];
			force_valid_4_3_mid_3 = 1'b0;
			force_valid_4_4_bottom_2 = 1'b0;
			force_valid_4_4_mid_2 = 1'b0;
			force_valid_4_4_top_1 = 1'b0;
			force_valid_1_2_bottom_2 = 1'b0;
			force_valid_1_2_mid_3 = 1'b0;
			end
		BINARY_231:
			begin
			force_valid_4_4_bottom_2 = neighbor_force_valid_1[14];
			force_valid_4_3_mid_3 = 1'b0;
			force_valid_4_3_top_2 = 1'b0;
			force_valid_4_4_mid_2 = 1'b0;
			force_valid_4_4_top_1 = 1'b0;
			force_valid_1_2_bottom_2 = 1'b0;
			force_valid_1_2_mid_3 = 1'b0;
			end
		BINARY_232:
			begin
			force_valid_4_4_mid_2 = neighbor_force_valid_1[14];
			force_valid_4_3_mid_3 = 1'b0;
			force_valid_4_3_top_2 = 1'b0;
			force_valid_4_4_bottom_2 = 1'b0;
			force_valid_4_4_top_1 = 1'b0;
			force_valid_1_2_bottom_2 = 1'b0;
			force_valid_1_2_mid_3 = 1'b0;
			end
		BINARY_233:
			begin
			force_valid_4_4_top_1 = neighbor_force_valid_1[14];
			force_valid_4_3_mid_3 = 1'b0;
			force_valid_4_3_top_2 = 1'b0;
			force_valid_4_4_bottom_2 = 1'b0;
			force_valid_4_4_mid_2 = 1'b0;
			force_valid_1_2_bottom_2 = 1'b0;
			force_valid_1_2_mid_3 = 1'b0;
			end
		BINARY_311:
			begin
			force_valid_1_2_bottom_2 = neighbor_force_valid_1[14];
			force_valid_4_3_mid_3 = 1'b0;
			force_valid_4_3_top_2 = 1'b0;
			force_valid_4_4_bottom_2 = 1'b0;
			force_valid_4_4_mid_2 = 1'b0;
			force_valid_4_4_top_1 = 1'b0;
			force_valid_1_2_mid_3 = 1'b0;
			end
		BINARY_312:
			begin
			force_valid_1_2_mid_3 = neighbor_force_valid_1[14];
			force_valid_4_3_mid_3 = 1'b0;
			force_valid_4_3_top_2 = 1'b0;
			force_valid_4_4_bottom_2 = 1'b0;
			force_valid_4_4_mid_2 = 1'b0;
			force_valid_4_4_top_1 = 1'b0;
			force_valid_1_2_bottom_2 = 1'b0;
			end
		default:
			begin
			force_valid_4_3_mid_3 = 1'b0;
			force_valid_4_3_top_2 = 1'b0;
			force_valid_4_4_bottom_2 = 1'b0;
			force_valid_4_4_mid_2 = 1'b0;
			force_valid_4_4_top_1 = 1'b0;
			force_valid_1_2_bottom_2 = 1'b0;
			force_valid_1_2_mid_3 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_1[15*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:15*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_222:
			begin
			force_valid_4_4_mid_3 = neighbor_force_valid_1[15];
			force_valid_4_4_top_2 = 1'b0;
			force_valid_4_1_bottom_2 = 1'b0;
			force_valid_4_1_mid_3 = 1'b0;
			force_valid_4_1_top_2 = 1'b0;
			force_valid_1_3_bottom_2 = 1'b0;
			force_valid_1_3_mid_3 = 1'b0;
			end
		BINARY_223:
			begin
			force_valid_4_4_top_2 = neighbor_force_valid_1[15];
			force_valid_4_4_mid_3 = 1'b0;
			force_valid_4_1_bottom_2 = 1'b0;
			force_valid_4_1_mid_3 = 1'b0;
			force_valid_4_1_top_2 = 1'b0;
			force_valid_1_3_bottom_2 = 1'b0;
			force_valid_1_3_mid_3 = 1'b0;
			end
		BINARY_231:
			begin
			force_valid_4_1_bottom_2 = neighbor_force_valid_1[15];
			force_valid_4_4_mid_3 = 1'b0;
			force_valid_4_4_top_2 = 1'b0;
			force_valid_4_1_mid_3 = 1'b0;
			force_valid_4_1_top_2 = 1'b0;
			force_valid_1_3_bottom_2 = 1'b0;
			force_valid_1_3_mid_3 = 1'b0;
			end
		BINARY_232:
			begin
			force_valid_4_1_mid_3 = neighbor_force_valid_1[15];
			force_valid_4_4_mid_3 = 1'b0;
			force_valid_4_4_top_2 = 1'b0;
			force_valid_4_1_bottom_2 = 1'b0;
			force_valid_4_1_top_2 = 1'b0;
			force_valid_1_3_bottom_2 = 1'b0;
			force_valid_1_3_mid_3 = 1'b0;
			end
		BINARY_233:
			begin
			force_valid_4_1_top_2 = neighbor_force_valid_1[15];
			force_valid_4_4_mid_3 = 1'b0;
			force_valid_4_4_top_2 = 1'b0;
			force_valid_4_1_bottom_2 = 1'b0;
			force_valid_4_1_mid_3 = 1'b0;
			force_valid_1_3_bottom_2 = 1'b0;
			force_valid_1_3_mid_3 = 1'b0;
			end
		BINARY_311:
			begin
			force_valid_1_3_bottom_2 = neighbor_force_valid_1[15];
			force_valid_4_4_mid_3 = 1'b0;
			force_valid_4_4_top_2 = 1'b0;
			force_valid_4_1_bottom_2 = 1'b0;
			force_valid_4_1_mid_3 = 1'b0;
			force_valid_4_1_top_2 = 1'b0;
			force_valid_1_3_mid_3 = 1'b0;
			end
		BINARY_312:
			begin
			force_valid_1_3_mid_3 = neighbor_force_valid_1[15];
			force_valid_4_4_mid_3 = 1'b0;
			force_valid_4_4_top_2 = 1'b0;
			force_valid_4_1_bottom_2 = 1'b0;
			force_valid_4_1_mid_3 = 1'b0;
			force_valid_4_1_top_2 = 1'b0;
			force_valid_1_3_bottom_2 = 1'b0;
			end
		default:
			begin
			force_valid_4_4_mid_3 = 1'b0;
			force_valid_4_4_top_2 = 1'b0;
			force_valid_4_1_bottom_2 = 1'b0;
			force_valid_4_1_mid_3 = 1'b0;
			force_valid_4_1_top_2 = 1'b0;
			force_valid_1_3_bottom_2 = 1'b0;
			force_valid_1_3_mid_3 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_2[0*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:0*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_313:
			begin
			force_valid_2_4_top_3 = neighbor_force_valid_2[0];
			force_valid_2_1_bottom_3 = 1'b0;
			force_valid_2_1_mid_4 = 1'b0;
			force_valid_2_1_top_3 = 1'b0;
			force_valid_2_2_bottom_3 = 1'b0;
			force_valid_2_2_mid_4 = 1'b0;
			force_valid_2_2_top_3 = 1'b0;
			end
		BINARY_321:
			begin
			force_valid_2_1_bottom_3 = neighbor_force_valid_2[0];
			force_valid_2_4_top_3 = 1'b0;
			force_valid_2_1_mid_4 = 1'b0;
			force_valid_2_1_top_3 = 1'b0;
			force_valid_2_2_bottom_3 = 1'b0;
			force_valid_2_2_mid_4 = 1'b0;
			force_valid_2_2_top_3 = 1'b0;
			end
		BINARY_322:
			begin
			force_valid_2_1_mid_4 = neighbor_force_valid_2[0];
			force_valid_2_4_top_3 = 1'b0;
			force_valid_2_1_bottom_3 = 1'b0;
			force_valid_2_1_top_3 = 1'b0;
			force_valid_2_2_bottom_3 = 1'b0;
			force_valid_2_2_mid_4 = 1'b0;
			force_valid_2_2_top_3 = 1'b0;
			end
		BINARY_323:
			begin
			force_valid_2_1_top_3 = neighbor_force_valid_2[0];
			force_valid_2_4_top_3 = 1'b0;
			force_valid_2_1_bottom_3 = 1'b0;
			force_valid_2_1_mid_4 = 1'b0;
			force_valid_2_2_bottom_3 = 1'b0;
			force_valid_2_2_mid_4 = 1'b0;
			force_valid_2_2_top_3 = 1'b0;
			end
		BINARY_331:
			begin
			force_valid_2_2_bottom_3 = neighbor_force_valid_2[0];
			force_valid_2_4_top_3 = 1'b0;
			force_valid_2_1_bottom_3 = 1'b0;
			force_valid_2_1_mid_4 = 1'b0;
			force_valid_2_1_top_3 = 1'b0;
			force_valid_2_2_mid_4 = 1'b0;
			force_valid_2_2_top_3 = 1'b0;
			end
		BINARY_332:
			begin
			force_valid_2_2_mid_4 = neighbor_force_valid_2[0];
			force_valid_2_4_top_3 = 1'b0;
			force_valid_2_1_bottom_3 = 1'b0;
			force_valid_2_1_mid_4 = 1'b0;
			force_valid_2_1_top_3 = 1'b0;
			force_valid_2_2_bottom_3 = 1'b0;
			force_valid_2_2_top_3 = 1'b0;
			end
		BINARY_333:
			begin
			force_valid_2_2_top_3 = neighbor_force_valid_2[0];
			force_valid_2_4_top_3 = 1'b0;
			force_valid_2_1_bottom_3 = 1'b0;
			force_valid_2_1_mid_4 = 1'b0;
			force_valid_2_1_top_3 = 1'b0;
			force_valid_2_2_bottom_3 = 1'b0;
			force_valid_2_2_mid_4 = 1'b0;
			end
		default:
			begin
			force_valid_2_4_top_3 = 1'b0;
			force_valid_2_1_bottom_3 = 1'b0;
			force_valid_2_1_mid_4 = 1'b0;
			force_valid_2_1_top_3 = 1'b0;
			force_valid_2_2_bottom_3 = 1'b0;
			force_valid_2_2_mid_4 = 1'b0;
			force_valid_2_2_top_3 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_2[1*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:1*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_313:
			begin
			force_valid_2_1_top_4 = neighbor_force_valid_2[1];
			force_valid_2_2_bottom_4 = 1'b0;
			force_valid_2_2_mid_5 = 1'b0;
			force_valid_2_2_top_4 = 1'b0;
			force_valid_2_3_bottom_3 = 1'b0;
			force_valid_2_3_mid_4 = 1'b0;
			force_valid_2_3_top_3 = 1'b0;
			end
		BINARY_321:
			begin
			force_valid_2_2_bottom_4 = neighbor_force_valid_2[1];
			force_valid_2_1_top_4 = 1'b0;
			force_valid_2_2_mid_5 = 1'b0;
			force_valid_2_2_top_4 = 1'b0;
			force_valid_2_3_bottom_3 = 1'b0;
			force_valid_2_3_mid_4 = 1'b0;
			force_valid_2_3_top_3 = 1'b0;
			end
		BINARY_322:
			begin
			force_valid_2_2_mid_5 = neighbor_force_valid_2[1];
			force_valid_2_1_top_4 = 1'b0;
			force_valid_2_2_bottom_4 = 1'b0;
			force_valid_2_2_top_4 = 1'b0;
			force_valid_2_3_bottom_3 = 1'b0;
			force_valid_2_3_mid_4 = 1'b0;
			force_valid_2_3_top_3 = 1'b0;
			end
		BINARY_323:
			begin
			force_valid_2_2_top_4 = neighbor_force_valid_2[1];
			force_valid_2_1_top_4 = 1'b0;
			force_valid_2_2_bottom_4 = 1'b0;
			force_valid_2_2_mid_5 = 1'b0;
			force_valid_2_3_bottom_3 = 1'b0;
			force_valid_2_3_mid_4 = 1'b0;
			force_valid_2_3_top_3 = 1'b0;
			end
		BINARY_331:
			begin
			force_valid_2_3_bottom_3 = neighbor_force_valid_2[1];
			force_valid_2_1_top_4 = 1'b0;
			force_valid_2_2_bottom_4 = 1'b0;
			force_valid_2_2_mid_5 = 1'b0;
			force_valid_2_2_top_4 = 1'b0;
			force_valid_2_3_mid_4 = 1'b0;
			force_valid_2_3_top_3 = 1'b0;
			end
		BINARY_332:
			begin
			force_valid_2_3_mid_4 = neighbor_force_valid_2[1];
			force_valid_2_1_top_4 = 1'b0;
			force_valid_2_2_bottom_4 = 1'b0;
			force_valid_2_2_mid_5 = 1'b0;
			force_valid_2_2_top_4 = 1'b0;
			force_valid_2_3_bottom_3 = 1'b0;
			force_valid_2_3_top_3 = 1'b0;
			end
		BINARY_333:
			begin
			force_valid_2_3_top_3 = neighbor_force_valid_2[1];
			force_valid_2_1_top_4 = 1'b0;
			force_valid_2_2_bottom_4 = 1'b0;
			force_valid_2_2_mid_5 = 1'b0;
			force_valid_2_2_top_4 = 1'b0;
			force_valid_2_3_bottom_3 = 1'b0;
			force_valid_2_3_mid_4 = 1'b0;
			end
		default:
			begin
			force_valid_2_1_top_4 = 1'b0;
			force_valid_2_2_bottom_4 = 1'b0;
			force_valid_2_2_mid_5 = 1'b0;
			force_valid_2_2_top_4 = 1'b0;
			force_valid_2_3_bottom_3 = 1'b0;
			force_valid_2_3_mid_4 = 1'b0;
			force_valid_2_3_top_3 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_2[2*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:2*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_313:
			begin
			force_valid_2_2_top_5 = neighbor_force_valid_2[2];
			force_valid_2_3_bottom_4 = 1'b0;
			force_valid_2_3_mid_5 = 1'b0;
			force_valid_2_3_top_4 = 1'b0;
			force_valid_2_4_bottom_3 = 1'b0;
			force_valid_2_4_mid_4 = 1'b0;
			force_valid_2_4_top_4 = 1'b0;
			end
		BINARY_321:
			begin
			force_valid_2_3_bottom_4 = neighbor_force_valid_2[2];
			force_valid_2_2_top_5 = 1'b0;
			force_valid_2_3_mid_5 = 1'b0;
			force_valid_2_3_top_4 = 1'b0;
			force_valid_2_4_bottom_3 = 1'b0;
			force_valid_2_4_mid_4 = 1'b0;
			force_valid_2_4_top_4 = 1'b0;
			end
		BINARY_322:
			begin
			force_valid_2_3_mid_5 = neighbor_force_valid_2[2];
			force_valid_2_2_top_5 = 1'b0;
			force_valid_2_3_bottom_4 = 1'b0;
			force_valid_2_3_top_4 = 1'b0;
			force_valid_2_4_bottom_3 = 1'b0;
			force_valid_2_4_mid_4 = 1'b0;
			force_valid_2_4_top_4 = 1'b0;
			end
		BINARY_323:
			begin
			force_valid_2_3_top_4 = neighbor_force_valid_2[2];
			force_valid_2_2_top_5 = 1'b0;
			force_valid_2_3_bottom_4 = 1'b0;
			force_valid_2_3_mid_5 = 1'b0;
			force_valid_2_4_bottom_3 = 1'b0;
			force_valid_2_4_mid_4 = 1'b0;
			force_valid_2_4_top_4 = 1'b0;
			end
		BINARY_331:
			begin
			force_valid_2_4_bottom_3 = neighbor_force_valid_2[2];
			force_valid_2_2_top_5 = 1'b0;
			force_valid_2_3_bottom_4 = 1'b0;
			force_valid_2_3_mid_5 = 1'b0;
			force_valid_2_3_top_4 = 1'b0;
			force_valid_2_4_mid_4 = 1'b0;
			force_valid_2_4_top_4 = 1'b0;
			end
		BINARY_332:
			begin
			force_valid_2_4_mid_4 = neighbor_force_valid_2[2];
			force_valid_2_2_top_5 = 1'b0;
			force_valid_2_3_bottom_4 = 1'b0;
			force_valid_2_3_mid_5 = 1'b0;
			force_valid_2_3_top_4 = 1'b0;
			force_valid_2_4_bottom_3 = 1'b0;
			force_valid_2_4_top_4 = 1'b0;
			end
		BINARY_333:
			begin
			force_valid_2_4_top_4 = neighbor_force_valid_2[2];
			force_valid_2_2_top_5 = 1'b0;
			force_valid_2_3_bottom_4 = 1'b0;
			force_valid_2_3_mid_5 = 1'b0;
			force_valid_2_3_top_4 = 1'b0;
			force_valid_2_4_bottom_3 = 1'b0;
			force_valid_2_4_mid_4 = 1'b0;
			end
		default:
			begin
			force_valid_2_2_top_5 = 1'b0;
			force_valid_2_3_bottom_4 = 1'b0;
			force_valid_2_3_mid_5 = 1'b0;
			force_valid_2_3_top_4 = 1'b0;
			force_valid_2_4_bottom_3 = 1'b0;
			force_valid_2_4_mid_4 = 1'b0;
			force_valid_2_4_top_4 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_2[3*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:3*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_313:
			begin
			force_valid_2_3_top_5 = neighbor_force_valid_2[3];
			force_valid_2_4_bottom_4 = 1'b0;
			force_valid_2_4_mid_5 = 1'b0;
			force_valid_2_4_top_5 = 1'b0;
			force_valid_2_1_bottom_4 = 1'b0;
			force_valid_2_1_mid_5 = 1'b0;
			force_valid_2_1_top_5 = 1'b0;
			end
		BINARY_321:
			begin
			force_valid_2_4_bottom_4 = neighbor_force_valid_2[3];
			force_valid_2_3_top_5 = 1'b0;
			force_valid_2_4_mid_5 = 1'b0;
			force_valid_2_4_top_5 = 1'b0;
			force_valid_2_1_bottom_4 = 1'b0;
			force_valid_2_1_mid_5 = 1'b0;
			force_valid_2_1_top_5 = 1'b0;
			end
		BINARY_322:
			begin
			force_valid_2_4_mid_5 = neighbor_force_valid_2[3];
			force_valid_2_3_top_5 = 1'b0;
			force_valid_2_4_bottom_4 = 1'b0;
			force_valid_2_4_top_5 = 1'b0;
			force_valid_2_1_bottom_4 = 1'b0;
			force_valid_2_1_mid_5 = 1'b0;
			force_valid_2_1_top_5 = 1'b0;
			end
		BINARY_323:
			begin
			force_valid_2_4_top_5 = neighbor_force_valid_2[3];
			force_valid_2_3_top_5 = 1'b0;
			force_valid_2_4_bottom_4 = 1'b0;
			force_valid_2_4_mid_5 = 1'b0;
			force_valid_2_1_bottom_4 = 1'b0;
			force_valid_2_1_mid_5 = 1'b0;
			force_valid_2_1_top_5 = 1'b0;
			end
		BINARY_331:
			begin
			force_valid_2_1_bottom_4 = neighbor_force_valid_2[3];
			force_valid_2_3_top_5 = 1'b0;
			force_valid_2_4_bottom_4 = 1'b0;
			force_valid_2_4_mid_5 = 1'b0;
			force_valid_2_4_top_5 = 1'b0;
			force_valid_2_1_mid_5 = 1'b0;
			force_valid_2_1_top_5 = 1'b0;
			end
		BINARY_332:
			begin
			force_valid_2_1_mid_5 = neighbor_force_valid_2[3];
			force_valid_2_3_top_5 = 1'b0;
			force_valid_2_4_bottom_4 = 1'b0;
			force_valid_2_4_mid_5 = 1'b0;
			force_valid_2_4_top_5 = 1'b0;
			force_valid_2_1_bottom_4 = 1'b0;
			force_valid_2_1_top_5 = 1'b0;
			end
		BINARY_333:
			begin
			force_valid_2_1_top_5 = neighbor_force_valid_2[3];
			force_valid_2_3_top_5 = 1'b0;
			force_valid_2_4_bottom_4 = 1'b0;
			force_valid_2_4_mid_5 = 1'b0;
			force_valid_2_4_top_5 = 1'b0;
			force_valid_2_1_bottom_4 = 1'b0;
			force_valid_2_1_mid_5 = 1'b0;
			end
		default:
			begin
			force_valid_2_3_top_5 = 1'b0;
			force_valid_2_4_bottom_4 = 1'b0;
			force_valid_2_4_mid_5 = 1'b0;
			force_valid_2_4_top_5 = 1'b0;
			force_valid_2_1_bottom_4 = 1'b0;
			force_valid_2_1_mid_5 = 1'b0;
			force_valid_2_1_top_5 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_2[4*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:4*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_313:
			begin
			force_valid_3_4_top_3 = neighbor_force_valid_2[4];
			force_valid_3_1_bottom_3 = 1'b0;
			force_valid_3_1_mid_4 = 1'b0;
			force_valid_3_1_top_3 = 1'b0;
			force_valid_3_2_bottom_3 = 1'b0;
			force_valid_3_2_mid_4 = 1'b0;
			force_valid_3_2_top_3 = 1'b0;
			end
		BINARY_321:
			begin
			force_valid_3_1_bottom_3 = neighbor_force_valid_2[4];
			force_valid_3_4_top_3 = 1'b0;
			force_valid_3_1_mid_4 = 1'b0;
			force_valid_3_1_top_3 = 1'b0;
			force_valid_3_2_bottom_3 = 1'b0;
			force_valid_3_2_mid_4 = 1'b0;
			force_valid_3_2_top_3 = 1'b0;
			end
		BINARY_322:
			begin
			force_valid_3_1_mid_4 = neighbor_force_valid_2[4];
			force_valid_3_4_top_3 = 1'b0;
			force_valid_3_1_bottom_3 = 1'b0;
			force_valid_3_1_top_3 = 1'b0;
			force_valid_3_2_bottom_3 = 1'b0;
			force_valid_3_2_mid_4 = 1'b0;
			force_valid_3_2_top_3 = 1'b0;
			end
		BINARY_323:
			begin
			force_valid_3_1_top_3 = neighbor_force_valid_2[4];
			force_valid_3_4_top_3 = 1'b0;
			force_valid_3_1_bottom_3 = 1'b0;
			force_valid_3_1_mid_4 = 1'b0;
			force_valid_3_2_bottom_3 = 1'b0;
			force_valid_3_2_mid_4 = 1'b0;
			force_valid_3_2_top_3 = 1'b0;
			end
		BINARY_331:
			begin
			force_valid_3_2_bottom_3 = neighbor_force_valid_2[4];
			force_valid_3_4_top_3 = 1'b0;
			force_valid_3_1_bottom_3 = 1'b0;
			force_valid_3_1_mid_4 = 1'b0;
			force_valid_3_1_top_3 = 1'b0;
			force_valid_3_2_mid_4 = 1'b0;
			force_valid_3_2_top_3 = 1'b0;
			end
		BINARY_332:
			begin
			force_valid_3_2_mid_4 = neighbor_force_valid_2[4];
			force_valid_3_4_top_3 = 1'b0;
			force_valid_3_1_bottom_3 = 1'b0;
			force_valid_3_1_mid_4 = 1'b0;
			force_valid_3_1_top_3 = 1'b0;
			force_valid_3_2_bottom_3 = 1'b0;
			force_valid_3_2_top_3 = 1'b0;
			end
		BINARY_333:
			begin
			force_valid_3_2_top_3 = neighbor_force_valid_2[4];
			force_valid_3_4_top_3 = 1'b0;
			force_valid_3_1_bottom_3 = 1'b0;
			force_valid_3_1_mid_4 = 1'b0;
			force_valid_3_1_top_3 = 1'b0;
			force_valid_3_2_bottom_3 = 1'b0;
			force_valid_3_2_mid_4 = 1'b0;
			end
		default:
			begin
			force_valid_3_4_top_3 = 1'b0;
			force_valid_3_1_bottom_3 = 1'b0;
			force_valid_3_1_mid_4 = 1'b0;
			force_valid_3_1_top_3 = 1'b0;
			force_valid_3_2_bottom_3 = 1'b0;
			force_valid_3_2_mid_4 = 1'b0;
			force_valid_3_2_top_3 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_2[5*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:5*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_313:
			begin
			force_valid_3_1_top_4 = neighbor_force_valid_2[5];
			force_valid_3_2_bottom_4 = 1'b0;
			force_valid_3_2_mid_5 = 1'b0;
			force_valid_3_2_top_4 = 1'b0;
			force_valid_3_3_bottom_3 = 1'b0;
			force_valid_3_3_mid_4 = 1'b0;
			force_valid_3_3_top_3 = 1'b0;
			end
		BINARY_321:
			begin
			force_valid_3_2_bottom_4 = neighbor_force_valid_2[5];
			force_valid_3_1_top_4 = 1'b0;
			force_valid_3_2_mid_5 = 1'b0;
			force_valid_3_2_top_4 = 1'b0;
			force_valid_3_3_bottom_3 = 1'b0;
			force_valid_3_3_mid_4 = 1'b0;
			force_valid_3_3_top_3 = 1'b0;
			end
		BINARY_322:
			begin
			force_valid_3_2_mid_5 = neighbor_force_valid_2[5];
			force_valid_3_1_top_4 = 1'b0;
			force_valid_3_2_bottom_4 = 1'b0;
			force_valid_3_2_top_4 = 1'b0;
			force_valid_3_3_bottom_3 = 1'b0;
			force_valid_3_3_mid_4 = 1'b0;
			force_valid_3_3_top_3 = 1'b0;
			end
		BINARY_323:
			begin
			force_valid_3_2_top_4 = neighbor_force_valid_2[5];
			force_valid_3_1_top_4 = 1'b0;
			force_valid_3_2_bottom_4 = 1'b0;
			force_valid_3_2_mid_5 = 1'b0;
			force_valid_3_3_bottom_3 = 1'b0;
			force_valid_3_3_mid_4 = 1'b0;
			force_valid_3_3_top_3 = 1'b0;
			end
		BINARY_331:
			begin
			force_valid_3_3_bottom_3 = neighbor_force_valid_2[5];
			force_valid_3_1_top_4 = 1'b0;
			force_valid_3_2_bottom_4 = 1'b0;
			force_valid_3_2_mid_5 = 1'b0;
			force_valid_3_2_top_4 = 1'b0;
			force_valid_3_3_mid_4 = 1'b0;
			force_valid_3_3_top_3 = 1'b0;
			end
		BINARY_332:
			begin
			force_valid_3_3_mid_4 = neighbor_force_valid_2[5];
			force_valid_3_1_top_4 = 1'b0;
			force_valid_3_2_bottom_4 = 1'b0;
			force_valid_3_2_mid_5 = 1'b0;
			force_valid_3_2_top_4 = 1'b0;
			force_valid_3_3_bottom_3 = 1'b0;
			force_valid_3_3_top_3 = 1'b0;
			end
		BINARY_333:
			begin
			force_valid_3_3_top_3 = neighbor_force_valid_2[5];
			force_valid_3_1_top_4 = 1'b0;
			force_valid_3_2_bottom_4 = 1'b0;
			force_valid_3_2_mid_5 = 1'b0;
			force_valid_3_2_top_4 = 1'b0;
			force_valid_3_3_bottom_3 = 1'b0;
			force_valid_3_3_mid_4 = 1'b0;
			end
		default:
			begin
			force_valid_3_1_top_4 = 1'b0;
			force_valid_3_2_bottom_4 = 1'b0;
			force_valid_3_2_mid_5 = 1'b0;
			force_valid_3_2_top_4 = 1'b0;
			force_valid_3_3_bottom_3 = 1'b0;
			force_valid_3_3_mid_4 = 1'b0;
			force_valid_3_3_top_3 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_2[6*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:6*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_313:
			begin
			force_valid_3_2_top_5 = neighbor_force_valid_2[6];
			force_valid_3_3_bottom_4 = 1'b0;
			force_valid_3_3_mid_5 = 1'b0;
			force_valid_3_3_top_4 = 1'b0;
			force_valid_3_4_bottom_3 = 1'b0;
			force_valid_3_4_mid_4 = 1'b0;
			force_valid_3_4_top_4 = 1'b0;
			end
		BINARY_321:
			begin
			force_valid_3_3_bottom_4 = neighbor_force_valid_2[6];
			force_valid_3_2_top_5 = 1'b0;
			force_valid_3_3_mid_5 = 1'b0;
			force_valid_3_3_top_4 = 1'b0;
			force_valid_3_4_bottom_3 = 1'b0;
			force_valid_3_4_mid_4 = 1'b0;
			force_valid_3_4_top_4 = 1'b0;
			end
		BINARY_322:
			begin
			force_valid_3_3_mid_5 = neighbor_force_valid_2[6];
			force_valid_3_2_top_5 = 1'b0;
			force_valid_3_3_bottom_4 = 1'b0;
			force_valid_3_3_top_4 = 1'b0;
			force_valid_3_4_bottom_3 = 1'b0;
			force_valid_3_4_mid_4 = 1'b0;
			force_valid_3_4_top_4 = 1'b0;
			end
		BINARY_323:
			begin
			force_valid_3_3_top_4 = neighbor_force_valid_2[6];
			force_valid_3_2_top_5 = 1'b0;
			force_valid_3_3_bottom_4 = 1'b0;
			force_valid_3_3_mid_5 = 1'b0;
			force_valid_3_4_bottom_3 = 1'b0;
			force_valid_3_4_mid_4 = 1'b0;
			force_valid_3_4_top_4 = 1'b0;
			end
		BINARY_331:
			begin
			force_valid_3_4_bottom_3 = neighbor_force_valid_2[6];
			force_valid_3_2_top_5 = 1'b0;
			force_valid_3_3_bottom_4 = 1'b0;
			force_valid_3_3_mid_5 = 1'b0;
			force_valid_3_3_top_4 = 1'b0;
			force_valid_3_4_mid_4 = 1'b0;
			force_valid_3_4_top_4 = 1'b0;
			end
		BINARY_332:
			begin
			force_valid_3_4_mid_4 = neighbor_force_valid_2[6];
			force_valid_3_2_top_5 = 1'b0;
			force_valid_3_3_bottom_4 = 1'b0;
			force_valid_3_3_mid_5 = 1'b0;
			force_valid_3_3_top_4 = 1'b0;
			force_valid_3_4_bottom_3 = 1'b0;
			force_valid_3_4_top_4 = 1'b0;
			end
		BINARY_333:
			begin
			force_valid_3_4_top_4 = neighbor_force_valid_2[6];
			force_valid_3_2_top_5 = 1'b0;
			force_valid_3_3_bottom_4 = 1'b0;
			force_valid_3_3_mid_5 = 1'b0;
			force_valid_3_3_top_4 = 1'b0;
			force_valid_3_4_bottom_3 = 1'b0;
			force_valid_3_4_mid_4 = 1'b0;
			end
		default:
			begin
			force_valid_3_2_top_5 = 1'b0;
			force_valid_3_3_bottom_4 = 1'b0;
			force_valid_3_3_mid_5 = 1'b0;
			force_valid_3_3_top_4 = 1'b0;
			force_valid_3_4_bottom_3 = 1'b0;
			force_valid_3_4_mid_4 = 1'b0;
			force_valid_3_4_top_4 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_2[7*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:7*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_313:
			begin
			force_valid_3_3_top_5 = neighbor_force_valid_2[7];
			force_valid_3_4_bottom_4 = 1'b0;
			force_valid_3_4_mid_5 = 1'b0;
			force_valid_3_4_top_5 = 1'b0;
			force_valid_3_1_bottom_4 = 1'b0;
			force_valid_3_1_mid_5 = 1'b0;
			force_valid_3_1_top_5 = 1'b0;
			end
		BINARY_321:
			begin
			force_valid_3_4_bottom_4 = neighbor_force_valid_2[7];
			force_valid_3_3_top_5 = 1'b0;
			force_valid_3_4_mid_5 = 1'b0;
			force_valid_3_4_top_5 = 1'b0;
			force_valid_3_1_bottom_4 = 1'b0;
			force_valid_3_1_mid_5 = 1'b0;
			force_valid_3_1_top_5 = 1'b0;
			end
		BINARY_322:
			begin
			force_valid_3_4_mid_5 = neighbor_force_valid_2[7];
			force_valid_3_3_top_5 = 1'b0;
			force_valid_3_4_bottom_4 = 1'b0;
			force_valid_3_4_top_5 = 1'b0;
			force_valid_3_1_bottom_4 = 1'b0;
			force_valid_3_1_mid_5 = 1'b0;
			force_valid_3_1_top_5 = 1'b0;
			end
		BINARY_323:
			begin
			force_valid_3_4_top_5 = neighbor_force_valid_2[7];
			force_valid_3_3_top_5 = 1'b0;
			force_valid_3_4_bottom_4 = 1'b0;
			force_valid_3_4_mid_5 = 1'b0;
			force_valid_3_1_bottom_4 = 1'b0;
			force_valid_3_1_mid_5 = 1'b0;
			force_valid_3_1_top_5 = 1'b0;
			end
		BINARY_331:
			begin
			force_valid_3_1_bottom_4 = neighbor_force_valid_2[7];
			force_valid_3_3_top_5 = 1'b0;
			force_valid_3_4_bottom_4 = 1'b0;
			force_valid_3_4_mid_5 = 1'b0;
			force_valid_3_4_top_5 = 1'b0;
			force_valid_3_1_mid_5 = 1'b0;
			force_valid_3_1_top_5 = 1'b0;
			end
		BINARY_332:
			begin
			force_valid_3_1_mid_5 = neighbor_force_valid_2[7];
			force_valid_3_3_top_5 = 1'b0;
			force_valid_3_4_bottom_4 = 1'b0;
			force_valid_3_4_mid_5 = 1'b0;
			force_valid_3_4_top_5 = 1'b0;
			force_valid_3_1_bottom_4 = 1'b0;
			force_valid_3_1_top_5 = 1'b0;
			end
		BINARY_333:
			begin
			force_valid_3_1_top_5 = neighbor_force_valid_2[7];
			force_valid_3_3_top_5 = 1'b0;
			force_valid_3_4_bottom_4 = 1'b0;
			force_valid_3_4_mid_5 = 1'b0;
			force_valid_3_4_top_5 = 1'b0;
			force_valid_3_1_bottom_4 = 1'b0;
			force_valid_3_1_mid_5 = 1'b0;
			end
		default:
			begin
			force_valid_3_3_top_5 = 1'b0;
			force_valid_3_4_bottom_4 = 1'b0;
			force_valid_3_4_mid_5 = 1'b0;
			force_valid_3_4_top_5 = 1'b0;
			force_valid_3_1_bottom_4 = 1'b0;
			force_valid_3_1_mid_5 = 1'b0;
			force_valid_3_1_top_5 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_2[8*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:8*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_313:
			begin
			force_valid_4_4_top_3 = neighbor_force_valid_2[8];
			force_valid_4_1_bottom_3 = 1'b0;
			force_valid_4_1_mid_4 = 1'b0;
			force_valid_4_1_top_3 = 1'b0;
			force_valid_4_2_bottom_3 = 1'b0;
			force_valid_4_2_mid_4 = 1'b0;
			force_valid_4_2_top_3 = 1'b0;
			end
		BINARY_321:
			begin
			force_valid_4_1_bottom_3 = neighbor_force_valid_2[8];
			force_valid_4_4_top_3 = 1'b0;
			force_valid_4_1_mid_4 = 1'b0;
			force_valid_4_1_top_3 = 1'b0;
			force_valid_4_2_bottom_3 = 1'b0;
			force_valid_4_2_mid_4 = 1'b0;
			force_valid_4_2_top_3 = 1'b0;
			end
		BINARY_322:
			begin
			force_valid_4_1_mid_4 = neighbor_force_valid_2[8];
			force_valid_4_4_top_3 = 1'b0;
			force_valid_4_1_bottom_3 = 1'b0;
			force_valid_4_1_top_3 = 1'b0;
			force_valid_4_2_bottom_3 = 1'b0;
			force_valid_4_2_mid_4 = 1'b0;
			force_valid_4_2_top_3 = 1'b0;
			end
		BINARY_323:
			begin
			force_valid_4_1_top_3 = neighbor_force_valid_2[8];
			force_valid_4_4_top_3 = 1'b0;
			force_valid_4_1_bottom_3 = 1'b0;
			force_valid_4_1_mid_4 = 1'b0;
			force_valid_4_2_bottom_3 = 1'b0;
			force_valid_4_2_mid_4 = 1'b0;
			force_valid_4_2_top_3 = 1'b0;
			end
		BINARY_331:
			begin
			force_valid_4_2_bottom_3 = neighbor_force_valid_2[8];
			force_valid_4_4_top_3 = 1'b0;
			force_valid_4_1_bottom_3 = 1'b0;
			force_valid_4_1_mid_4 = 1'b0;
			force_valid_4_1_top_3 = 1'b0;
			force_valid_4_2_mid_4 = 1'b0;
			force_valid_4_2_top_3 = 1'b0;
			end
		BINARY_332:
			begin
			force_valid_4_2_mid_4 = neighbor_force_valid_2[8];
			force_valid_4_4_top_3 = 1'b0;
			force_valid_4_1_bottom_3 = 1'b0;
			force_valid_4_1_mid_4 = 1'b0;
			force_valid_4_1_top_3 = 1'b0;
			force_valid_4_2_bottom_3 = 1'b0;
			force_valid_4_2_top_3 = 1'b0;
			end
		BINARY_333:
			begin
			force_valid_4_2_top_3 = neighbor_force_valid_2[8];
			force_valid_4_4_top_3 = 1'b0;
			force_valid_4_1_bottom_3 = 1'b0;
			force_valid_4_1_mid_4 = 1'b0;
			force_valid_4_1_top_3 = 1'b0;
			force_valid_4_2_bottom_3 = 1'b0;
			force_valid_4_2_mid_4 = 1'b0;
			end
		default:
			begin
			force_valid_4_4_top_3 = 1'b0;
			force_valid_4_1_bottom_3 = 1'b0;
			force_valid_4_1_mid_4 = 1'b0;
			force_valid_4_1_top_3 = 1'b0;
			force_valid_4_2_bottom_3 = 1'b0;
			force_valid_4_2_mid_4 = 1'b0;
			force_valid_4_2_top_3 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_2[9*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:9*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_313:
			begin
			force_valid_4_1_top_4 = neighbor_force_valid_2[9];
			force_valid_4_2_bottom_4 = 1'b0;
			force_valid_4_2_mid_5 = 1'b0;
			force_valid_4_2_top_4 = 1'b0;
			force_valid_4_3_bottom_3 = 1'b0;
			force_valid_4_3_mid_4 = 1'b0;
			force_valid_4_3_top_3 = 1'b0;
			end
		BINARY_321:
			begin
			force_valid_4_2_bottom_4 = neighbor_force_valid_2[9];
			force_valid_4_1_top_4 = 1'b0;
			force_valid_4_2_mid_5 = 1'b0;
			force_valid_4_2_top_4 = 1'b0;
			force_valid_4_3_bottom_3 = 1'b0;
			force_valid_4_3_mid_4 = 1'b0;
			force_valid_4_3_top_3 = 1'b0;
			end
		BINARY_322:
			begin
			force_valid_4_2_mid_5 = neighbor_force_valid_2[9];
			force_valid_4_1_top_4 = 1'b0;
			force_valid_4_2_bottom_4 = 1'b0;
			force_valid_4_2_top_4 = 1'b0;
			force_valid_4_3_bottom_3 = 1'b0;
			force_valid_4_3_mid_4 = 1'b0;
			force_valid_4_3_top_3 = 1'b0;
			end
		BINARY_323:
			begin
			force_valid_4_2_top_4 = neighbor_force_valid_2[9];
			force_valid_4_1_top_4 = 1'b0;
			force_valid_4_2_bottom_4 = 1'b0;
			force_valid_4_2_mid_5 = 1'b0;
			force_valid_4_3_bottom_3 = 1'b0;
			force_valid_4_3_mid_4 = 1'b0;
			force_valid_4_3_top_3 = 1'b0;
			end
		BINARY_331:
			begin
			force_valid_4_3_bottom_3 = neighbor_force_valid_2[9];
			force_valid_4_1_top_4 = 1'b0;
			force_valid_4_2_bottom_4 = 1'b0;
			force_valid_4_2_mid_5 = 1'b0;
			force_valid_4_2_top_4 = 1'b0;
			force_valid_4_3_mid_4 = 1'b0;
			force_valid_4_3_top_3 = 1'b0;
			end
		BINARY_332:
			begin
			force_valid_4_3_mid_4 = neighbor_force_valid_2[9];
			force_valid_4_1_top_4 = 1'b0;
			force_valid_4_2_bottom_4 = 1'b0;
			force_valid_4_2_mid_5 = 1'b0;
			force_valid_4_2_top_4 = 1'b0;
			force_valid_4_3_bottom_3 = 1'b0;
			force_valid_4_3_top_3 = 1'b0;
			end
		BINARY_333:
			begin
			force_valid_4_3_top_3 = neighbor_force_valid_2[9];
			force_valid_4_1_top_4 = 1'b0;
			force_valid_4_2_bottom_4 = 1'b0;
			force_valid_4_2_mid_5 = 1'b0;
			force_valid_4_2_top_4 = 1'b0;
			force_valid_4_3_bottom_3 = 1'b0;
			force_valid_4_3_mid_4 = 1'b0;
			end
		default:
			begin
			force_valid_4_1_top_4 = 1'b0;
			force_valid_4_2_bottom_4 = 1'b0;
			force_valid_4_2_mid_5 = 1'b0;
			force_valid_4_2_top_4 = 1'b0;
			force_valid_4_3_bottom_3 = 1'b0;
			force_valid_4_3_mid_4 = 1'b0;
			force_valid_4_3_top_3 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_2[10*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:10*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_313:
			begin
			force_valid_4_2_top_5 = neighbor_force_valid_2[10];
			force_valid_4_3_bottom_4 = 1'b0;
			force_valid_4_3_mid_5 = 1'b0;
			force_valid_4_3_top_4 = 1'b0;
			force_valid_4_4_bottom_3 = 1'b0;
			force_valid_4_4_mid_4 = 1'b0;
			force_valid_4_4_top_4 = 1'b0;
			end
		BINARY_321:
			begin
			force_valid_4_3_bottom_4 = neighbor_force_valid_2[10];
			force_valid_4_2_top_5 = 1'b0;
			force_valid_4_3_mid_5 = 1'b0;
			force_valid_4_3_top_4 = 1'b0;
			force_valid_4_4_bottom_3 = 1'b0;
			force_valid_4_4_mid_4 = 1'b0;
			force_valid_4_4_top_4 = 1'b0;
			end
		BINARY_322:
			begin
			force_valid_4_3_mid_5 = neighbor_force_valid_2[10];
			force_valid_4_2_top_5 = 1'b0;
			force_valid_4_3_bottom_4 = 1'b0;
			force_valid_4_3_top_4 = 1'b0;
			force_valid_4_4_bottom_3 = 1'b0;
			force_valid_4_4_mid_4 = 1'b0;
			force_valid_4_4_top_4 = 1'b0;
			end
		BINARY_323:
			begin
			force_valid_4_3_top_4 = neighbor_force_valid_2[10];
			force_valid_4_2_top_5 = 1'b0;
			force_valid_4_3_bottom_4 = 1'b0;
			force_valid_4_3_mid_5 = 1'b0;
			force_valid_4_4_bottom_3 = 1'b0;
			force_valid_4_4_mid_4 = 1'b0;
			force_valid_4_4_top_4 = 1'b0;
			end
		BINARY_331:
			begin
			force_valid_4_4_bottom_3 = neighbor_force_valid_2[10];
			force_valid_4_2_top_5 = 1'b0;
			force_valid_4_3_bottom_4 = 1'b0;
			force_valid_4_3_mid_5 = 1'b0;
			force_valid_4_3_top_4 = 1'b0;
			force_valid_4_4_mid_4 = 1'b0;
			force_valid_4_4_top_4 = 1'b0;
			end
		BINARY_332:
			begin
			force_valid_4_4_mid_4 = neighbor_force_valid_2[10];
			force_valid_4_2_top_5 = 1'b0;
			force_valid_4_3_bottom_4 = 1'b0;
			force_valid_4_3_mid_5 = 1'b0;
			force_valid_4_3_top_4 = 1'b0;
			force_valid_4_4_bottom_3 = 1'b0;
			force_valid_4_4_top_4 = 1'b0;
			end
		BINARY_333:
			begin
			force_valid_4_4_top_4 = neighbor_force_valid_2[10];
			force_valid_4_2_top_5 = 1'b0;
			force_valid_4_3_bottom_4 = 1'b0;
			force_valid_4_3_mid_5 = 1'b0;
			force_valid_4_3_top_4 = 1'b0;
			force_valid_4_4_bottom_3 = 1'b0;
			force_valid_4_4_mid_4 = 1'b0;
			end
		default:
			begin
			force_valid_4_2_top_5 = 1'b0;
			force_valid_4_3_bottom_4 = 1'b0;
			force_valid_4_3_mid_5 = 1'b0;
			force_valid_4_3_top_4 = 1'b0;
			force_valid_4_4_bottom_3 = 1'b0;
			force_valid_4_4_mid_4 = 1'b0;
			force_valid_4_4_top_4 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_2[11*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:11*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_313:
			begin
			force_valid_4_3_top_5 = neighbor_force_valid_2[11];
			force_valid_4_4_bottom_4 = 1'b0;
			force_valid_4_4_mid_5 = 1'b0;
			force_valid_4_4_top_5 = 1'b0;
			force_valid_4_1_bottom_4 = 1'b0;
			force_valid_4_1_mid_5 = 1'b0;
			force_valid_4_1_top_5 = 1'b0;
			end
		BINARY_321:
			begin
			force_valid_4_4_bottom_4 = neighbor_force_valid_2[11];
			force_valid_4_3_top_5 = 1'b0;
			force_valid_4_4_mid_5 = 1'b0;
			force_valid_4_4_top_5 = 1'b0;
			force_valid_4_1_bottom_4 = 1'b0;
			force_valid_4_1_mid_5 = 1'b0;
			force_valid_4_1_top_5 = 1'b0;
			end
		BINARY_322:
			begin
			force_valid_4_4_mid_5 = neighbor_force_valid_2[11];
			force_valid_4_3_top_5 = 1'b0;
			force_valid_4_4_bottom_4 = 1'b0;
			force_valid_4_4_top_5 = 1'b0;
			force_valid_4_1_bottom_4 = 1'b0;
			force_valid_4_1_mid_5 = 1'b0;
			force_valid_4_1_top_5 = 1'b0;
			end
		BINARY_323:
			begin
			force_valid_4_4_top_5 = neighbor_force_valid_2[11];
			force_valid_4_3_top_5 = 1'b0;
			force_valid_4_4_bottom_4 = 1'b0;
			force_valid_4_4_mid_5 = 1'b0;
			force_valid_4_1_bottom_4 = 1'b0;
			force_valid_4_1_mid_5 = 1'b0;
			force_valid_4_1_top_5 = 1'b0;
			end
		BINARY_331:
			begin
			force_valid_4_1_bottom_4 = neighbor_force_valid_2[11];
			force_valid_4_3_top_5 = 1'b0;
			force_valid_4_4_bottom_4 = 1'b0;
			force_valid_4_4_mid_5 = 1'b0;
			force_valid_4_4_top_5 = 1'b0;
			force_valid_4_1_mid_5 = 1'b0;
			force_valid_4_1_top_5 = 1'b0;
			end
		BINARY_332:
			begin
			force_valid_4_1_mid_5 = neighbor_force_valid_2[11];
			force_valid_4_3_top_5 = 1'b0;
			force_valid_4_4_bottom_4 = 1'b0;
			force_valid_4_4_mid_5 = 1'b0;
			force_valid_4_4_top_5 = 1'b0;
			force_valid_4_1_bottom_4 = 1'b0;
			force_valid_4_1_top_5 = 1'b0;
			end
		BINARY_333:
			begin
			force_valid_4_1_top_5 = neighbor_force_valid_2[11];
			force_valid_4_3_top_5 = 1'b0;
			force_valid_4_4_bottom_4 = 1'b0;
			force_valid_4_4_mid_5 = 1'b0;
			force_valid_4_4_top_5 = 1'b0;
			force_valid_4_1_bottom_4 = 1'b0;
			force_valid_4_1_mid_5 = 1'b0;
			end
		default:
			begin
			force_valid_4_3_top_5 = 1'b0;
			force_valid_4_4_bottom_4 = 1'b0;
			force_valid_4_4_mid_5 = 1'b0;
			force_valid_4_4_top_5 = 1'b0;
			force_valid_4_1_bottom_4 = 1'b0;
			force_valid_4_1_mid_5 = 1'b0;
			force_valid_4_1_top_5 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_2[12*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:12*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_313:
			begin
			force_valid_1_4_top_3 = neighbor_force_valid_2[12];
			force_valid_1_1_bottom_3 = 1'b0;
			force_valid_1_1_mid_4 = 1'b0;
			force_valid_1_1_top_3 = 1'b0;
			force_valid_1_2_bottom_3 = 1'b0;
			force_valid_1_2_mid_4 = 1'b0;
			force_valid_1_2_top_3 = 1'b0;
			end
		BINARY_321:
			begin
			force_valid_1_1_bottom_3 = neighbor_force_valid_2[12];
			force_valid_1_4_top_3 = 1'b0;
			force_valid_1_1_mid_4 = 1'b0;
			force_valid_1_1_top_3 = 1'b0;
			force_valid_1_2_bottom_3 = 1'b0;
			force_valid_1_2_mid_4 = 1'b0;
			force_valid_1_2_top_3 = 1'b0;
			end
		BINARY_322:
			begin
			force_valid_1_1_mid_4 = neighbor_force_valid_2[12];
			force_valid_1_4_top_3 = 1'b0;
			force_valid_1_1_bottom_3 = 1'b0;
			force_valid_1_1_top_3 = 1'b0;
			force_valid_1_2_bottom_3 = 1'b0;
			force_valid_1_2_mid_4 = 1'b0;
			force_valid_1_2_top_3 = 1'b0;
			end
		BINARY_323:
			begin
			force_valid_1_1_top_3 = neighbor_force_valid_2[12];
			force_valid_1_4_top_3 = 1'b0;
			force_valid_1_1_bottom_3 = 1'b0;
			force_valid_1_1_mid_4 = 1'b0;
			force_valid_1_2_bottom_3 = 1'b0;
			force_valid_1_2_mid_4 = 1'b0;
			force_valid_1_2_top_3 = 1'b0;
			end
		BINARY_331:
			begin
			force_valid_1_2_bottom_3 = neighbor_force_valid_2[12];
			force_valid_1_4_top_3 = 1'b0;
			force_valid_1_1_bottom_3 = 1'b0;
			force_valid_1_1_mid_4 = 1'b0;
			force_valid_1_1_top_3 = 1'b0;
			force_valid_1_2_mid_4 = 1'b0;
			force_valid_1_2_top_3 = 1'b0;
			end
		BINARY_332:
			begin
			force_valid_1_2_mid_4 = neighbor_force_valid_2[12];
			force_valid_1_4_top_3 = 1'b0;
			force_valid_1_1_bottom_3 = 1'b0;
			force_valid_1_1_mid_4 = 1'b0;
			force_valid_1_1_top_3 = 1'b0;
			force_valid_1_2_bottom_3 = 1'b0;
			force_valid_1_2_top_3 = 1'b0;
			end
		BINARY_333:
			begin
			force_valid_1_2_top_3 = neighbor_force_valid_2[12];
			force_valid_1_4_top_3 = 1'b0;
			force_valid_1_1_bottom_3 = 1'b0;
			force_valid_1_1_mid_4 = 1'b0;
			force_valid_1_1_top_3 = 1'b0;
			force_valid_1_2_bottom_3 = 1'b0;
			force_valid_1_2_mid_4 = 1'b0;
			end
		default:
			begin
			force_valid_1_4_top_3 = 1'b0;
			force_valid_1_1_bottom_3 = 1'b0;
			force_valid_1_1_mid_4 = 1'b0;
			force_valid_1_1_top_3 = 1'b0;
			force_valid_1_2_bottom_3 = 1'b0;
			force_valid_1_2_mid_4 = 1'b0;
			force_valid_1_2_top_3 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_2[13*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:13*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_313:
			begin
			force_valid_1_1_top_4 = neighbor_force_valid_2[13];
			force_valid_1_2_bottom_4 = 1'b0;
			force_valid_1_2_mid_5 = 1'b0;
			force_valid_1_2_top_4 = 1'b0;
			force_valid_1_3_bottom_3 = 1'b0;
			force_valid_1_3_mid_4 = 1'b0;
			force_valid_1_3_top_3 = 1'b0;
			end
		BINARY_321:
			begin
			force_valid_1_2_bottom_4 = neighbor_force_valid_2[13];
			force_valid_1_1_top_4 = 1'b0;
			force_valid_1_2_mid_5 = 1'b0;
			force_valid_1_2_top_4 = 1'b0;
			force_valid_1_3_bottom_3 = 1'b0;
			force_valid_1_3_mid_4 = 1'b0;
			force_valid_1_3_top_3 = 1'b0;
			end
		BINARY_322:
			begin
			force_valid_1_2_mid_5 = neighbor_force_valid_2[13];
			force_valid_1_1_top_4 = 1'b0;
			force_valid_1_2_bottom_4 = 1'b0;
			force_valid_1_2_top_4 = 1'b0;
			force_valid_1_3_bottom_3 = 1'b0;
			force_valid_1_3_mid_4 = 1'b0;
			force_valid_1_3_top_3 = 1'b0;
			end
		BINARY_323:
			begin
			force_valid_1_2_top_4 = neighbor_force_valid_2[13];
			force_valid_1_1_top_4 = 1'b0;
			force_valid_1_2_bottom_4 = 1'b0;
			force_valid_1_2_mid_5 = 1'b0;
			force_valid_1_3_bottom_3 = 1'b0;
			force_valid_1_3_mid_4 = 1'b0;
			force_valid_1_3_top_3 = 1'b0;
			end
		BINARY_331:
			begin
			force_valid_1_3_bottom_3 = neighbor_force_valid_2[13];
			force_valid_1_1_top_4 = 1'b0;
			force_valid_1_2_bottom_4 = 1'b0;
			force_valid_1_2_mid_5 = 1'b0;
			force_valid_1_2_top_4 = 1'b0;
			force_valid_1_3_mid_4 = 1'b0;
			force_valid_1_3_top_3 = 1'b0;
			end
		BINARY_332:
			begin
			force_valid_1_3_mid_4 = neighbor_force_valid_2[13];
			force_valid_1_1_top_4 = 1'b0;
			force_valid_1_2_bottom_4 = 1'b0;
			force_valid_1_2_mid_5 = 1'b0;
			force_valid_1_2_top_4 = 1'b0;
			force_valid_1_3_bottom_3 = 1'b0;
			force_valid_1_3_top_3 = 1'b0;
			end
		BINARY_333:
			begin
			force_valid_1_3_top_3 = neighbor_force_valid_2[13];
			force_valid_1_1_top_4 = 1'b0;
			force_valid_1_2_bottom_4 = 1'b0;
			force_valid_1_2_mid_5 = 1'b0;
			force_valid_1_2_top_4 = 1'b0;
			force_valid_1_3_bottom_3 = 1'b0;
			force_valid_1_3_mid_4 = 1'b0;
			end
		default:
			begin
			force_valid_1_1_top_4 = 1'b0;
			force_valid_1_2_bottom_4 = 1'b0;
			force_valid_1_2_mid_5 = 1'b0;
			force_valid_1_2_top_4 = 1'b0;
			force_valid_1_3_bottom_3 = 1'b0;
			force_valid_1_3_mid_4 = 1'b0;
			force_valid_1_3_top_3 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_2[14*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:14*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_313:
			begin
			force_valid_1_2_top_5 = neighbor_force_valid_2[14];
			force_valid_1_3_bottom_4 = 1'b0;
			force_valid_1_3_mid_5 = 1'b0;
			force_valid_1_3_top_4 = 1'b0;
			force_valid_1_4_bottom_3 = 1'b0;
			force_valid_1_4_mid_4 = 1'b0;
			force_valid_1_4_top_4 = 1'b0;
			end
		BINARY_321:
			begin
			force_valid_1_3_bottom_4 = neighbor_force_valid_2[14];
			force_valid_1_2_top_5 = 1'b0;
			force_valid_1_3_mid_5 = 1'b0;
			force_valid_1_3_top_4 = 1'b0;
			force_valid_1_4_bottom_3 = 1'b0;
			force_valid_1_4_mid_4 = 1'b0;
			force_valid_1_4_top_4 = 1'b0;
			end
		BINARY_322:
			begin
			force_valid_1_3_mid_5 = neighbor_force_valid_2[14];
			force_valid_1_2_top_5 = 1'b0;
			force_valid_1_3_bottom_4 = 1'b0;
			force_valid_1_3_top_4 = 1'b0;
			force_valid_1_4_bottom_3 = 1'b0;
			force_valid_1_4_mid_4 = 1'b0;
			force_valid_1_4_top_4 = 1'b0;
			end
		BINARY_323:
			begin
			force_valid_1_3_top_4 = neighbor_force_valid_2[14];
			force_valid_1_2_top_5 = 1'b0;
			force_valid_1_3_bottom_4 = 1'b0;
			force_valid_1_3_mid_5 = 1'b0;
			force_valid_1_4_bottom_3 = 1'b0;
			force_valid_1_4_mid_4 = 1'b0;
			force_valid_1_4_top_4 = 1'b0;
			end
		BINARY_331:
			begin
			force_valid_1_4_bottom_3 = neighbor_force_valid_2[14];
			force_valid_1_2_top_5 = 1'b0;
			force_valid_1_3_bottom_4 = 1'b0;
			force_valid_1_3_mid_5 = 1'b0;
			force_valid_1_3_top_4 = 1'b0;
			force_valid_1_4_mid_4 = 1'b0;
			force_valid_1_4_top_4 = 1'b0;
			end
		BINARY_332:
			begin
			force_valid_1_4_mid_4 = neighbor_force_valid_2[14];
			force_valid_1_2_top_5 = 1'b0;
			force_valid_1_3_bottom_4 = 1'b0;
			force_valid_1_3_mid_5 = 1'b0;
			force_valid_1_3_top_4 = 1'b0;
			force_valid_1_4_bottom_3 = 1'b0;
			force_valid_1_4_top_4 = 1'b0;
			end
		BINARY_333:
			begin
			force_valid_1_4_top_4 = neighbor_force_valid_2[14];
			force_valid_1_2_top_5 = 1'b0;
			force_valid_1_3_bottom_4 = 1'b0;
			force_valid_1_3_mid_5 = 1'b0;
			force_valid_1_3_top_4 = 1'b0;
			force_valid_1_4_bottom_3 = 1'b0;
			force_valid_1_4_mid_4 = 1'b0;
			end
		default:
			begin
			force_valid_1_2_top_5 = 1'b0;
			force_valid_1_3_bottom_4 = 1'b0;
			force_valid_1_3_mid_5 = 1'b0;
			force_valid_1_3_top_4 = 1'b0;
			force_valid_1_4_bottom_3 = 1'b0;
			force_valid_1_4_mid_4 = 1'b0;
			force_valid_1_4_top_4 = 1'b0;
			end
	endcase
	end
always@(*)
	begin
	case(neighbor_force_data_from_FIFO_2[15*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH:15*FORCE_EVAL_FIFO_DATA_WIDTH+CELL_ADDR_WIDTH+1])
		BINARY_313:
			begin
			force_valid_1_3_top_5 = neighbor_force_valid_2[15];
			force_valid_1_4_bottom_4 = 1'b0;
			force_valid_1_4_mid_5 = 1'b0;
			force_valid_1_4_top_5 = 1'b0;
			force_valid_1_1_bottom_4 = 1'b0;
			force_valid_1_1_mid_5 = 1'b0;
			force_valid_1_1_top_5 = 1'b0;
			end
		BINARY_321:
			begin
			force_valid_1_4_bottom_4 = neighbor_force_valid_2[15];
			force_valid_1_3_top_5 = 1'b0;
			force_valid_1_4_mid_5 = 1'b0;
			force_valid_1_4_top_5 = 1'b0;
			force_valid_1_1_bottom_4 = 1'b0;
			force_valid_1_1_mid_5 = 1'b0;
			force_valid_1_1_top_5 = 1'b0;
			end
		BINARY_322:
			begin
			force_valid_1_4_mid_5 = neighbor_force_valid_2[15];
			force_valid_1_3_top_5 = 1'b0;
			force_valid_1_4_bottom_4 = 1'b0;
			force_valid_1_4_top_5 = 1'b0;
			force_valid_1_1_bottom_4 = 1'b0;
			force_valid_1_1_mid_5 = 1'b0;
			force_valid_1_1_top_5 = 1'b0;
			end
		BINARY_323:
			begin
			force_valid_1_4_top_5 = neighbor_force_valid_2[15];
			force_valid_1_3_top_5 = 1'b0;
			force_valid_1_4_bottom_4 = 1'b0;
			force_valid_1_4_mid_5 = 1'b0;
			force_valid_1_1_bottom_4 = 1'b0;
			force_valid_1_1_mid_5 = 1'b0;
			force_valid_1_1_top_5 = 1'b0;
			end
		BINARY_331:
			begin
			force_valid_1_1_bottom_4 = neighbor_force_valid_2[15];
			force_valid_1_3_top_5 = 1'b0;
			force_valid_1_4_bottom_4 = 1'b0;
			force_valid_1_4_mid_5 = 1'b0;
			force_valid_1_4_top_5 = 1'b0;
			force_valid_1_1_mid_5 = 1'b0;
			force_valid_1_1_top_5 = 1'b0;
			end
		BINARY_332:
			begin
			force_valid_1_1_mid_5 = neighbor_force_valid_2[15];
			force_valid_1_3_top_5 = 1'b0;
			force_valid_1_4_bottom_4 = 1'b0;
			force_valid_1_4_mid_5 = 1'b0;
			force_valid_1_4_top_5 = 1'b0;
			force_valid_1_1_bottom_4 = 1'b0;
			force_valid_1_1_top_5 = 1'b0;
			end
		BINARY_333:
			begin
			force_valid_1_1_top_5 = neighbor_force_valid_2[15];
			force_valid_1_3_top_5 = 1'b0;
			force_valid_1_4_bottom_4 = 1'b0;
			force_valid_1_4_mid_5 = 1'b0;
			force_valid_1_4_top_5 = 1'b0;
			force_valid_1_1_bottom_4 = 1'b0;
			force_valid_1_1_mid_5 = 1'b0;
			end
		default:
			begin
			force_valid_1_3_top_5 = 1'b0;
			force_valid_1_4_bottom_4 = 1'b0;
			force_valid_1_4_mid_5 = 1'b0;
			force_valid_1_4_top_5 = 1'b0;
			force_valid_1_1_bottom_4 = 1'b0;
			force_valid_1_1_mid_5 = 1'b0;
			force_valid_1_1_top_5 = 1'b0;
			end
	endcase
	end
	
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_1_1_mid
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(ref_force_valid[0]),
	.force_valid_1(force_valid_1_1_mid_1),
	.force_valid_2(force_valid_1_1_mid_2),
	.force_valid_3(force_valid_1_1_mid_3),
	.force_valid_4(force_valid_1_1_mid_4),
	.force_valid_5(force_valid_1_1_mid_5),

	.Arbitration_Result(Arbitration_1_1_mid)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_1_1_top
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_1_1_top_1),
	.force_valid_2(force_valid_1_1_top_2),
	.force_valid_3(force_valid_1_1_top_3),
	.force_valid_4(force_valid_1_1_top_4),
	.force_valid_5(force_valid_1_1_top_5),

	.Arbitration_Result(Arbitration_1_1_top)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_1_1_bottom
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_1_1_bottom_1),
	.force_valid_2(force_valid_1_1_bottom_2),
	.force_valid_3(force_valid_1_1_bottom_3),
	.force_valid_4(force_valid_1_1_bottom_4),
	.force_valid_5(1'b0),

	.Arbitration_Result(Arbitration_1_1_bottom)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_1_2_mid
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(ref_force_valid[1]),
	.force_valid_1(force_valid_1_2_mid_1),
	.force_valid_2(force_valid_1_2_mid_2),
	.force_valid_3(force_valid_1_2_mid_3),
	.force_valid_4(force_valid_1_2_mid_4),
	.force_valid_5(force_valid_1_2_mid_5),

	.Arbitration_Result(Arbitration_1_2_mid)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_1_2_top
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_1_2_top_1),
	.force_valid_2(force_valid_1_2_top_2),
	.force_valid_3(force_valid_1_2_top_3),
	.force_valid_4(force_valid_1_2_top_4),
	.force_valid_5(force_valid_1_2_top_5),

	.Arbitration_Result(Arbitration_1_2_top)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_1_2_bottom
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_1_2_bottom_1),
	.force_valid_2(force_valid_1_2_bottom_2),
	.force_valid_3(force_valid_1_2_bottom_3),
	.force_valid_4(force_valid_1_2_bottom_4),
	.force_valid_5(1'b0),

	.Arbitration_Result(Arbitration_1_2_bottom)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_1_3_mid
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(ref_force_valid[2]),
	.force_valid_1(force_valid_1_3_mid_1),
	.force_valid_2(force_valid_1_3_mid_2),
	.force_valid_3(force_valid_1_3_mid_3),
	.force_valid_4(force_valid_1_3_mid_4),
	.force_valid_5(force_valid_1_3_mid_5),

	.Arbitration_Result(Arbitration_1_3_mid)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_1_3_top
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_1_3_top_1),
	.force_valid_2(force_valid_1_3_top_2),
	.force_valid_3(force_valid_1_3_top_3),
	.force_valid_4(force_valid_1_3_top_4),
	.force_valid_5(force_valid_1_3_top_5),

	.Arbitration_Result(Arbitration_1_3_top)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_1_3_bottom
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_1_3_bottom_1),
	.force_valid_2(force_valid_1_3_bottom_2),
	.force_valid_3(force_valid_1_3_bottom_3),
	.force_valid_4(force_valid_1_3_bottom_4),
	.force_valid_5(1'b0),

	.Arbitration_Result(Arbitration_1_3_bottom)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_1_4_mid
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(ref_force_valid[3]),
	.force_valid_1(force_valid_1_4_mid_1),
	.force_valid_2(force_valid_1_4_mid_2),
	.force_valid_3(force_valid_1_4_mid_3),
	.force_valid_4(force_valid_1_4_mid_4),
	.force_valid_5(force_valid_1_4_mid_5),

	.Arbitration_Result(Arbitration_1_4_mid)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_1_4_top
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_1_4_top_1),
	.force_valid_2(force_valid_1_4_top_2),
	.force_valid_3(force_valid_1_4_top_3),
	.force_valid_4(force_valid_1_4_top_4),
	.force_valid_5(force_valid_1_4_top_5),

	.Arbitration_Result(Arbitration_1_4_top)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_1_4_bottom
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_1_4_bottom_1),
	.force_valid_2(force_valid_1_4_bottom_2),
	.force_valid_3(force_valid_1_4_bottom_3),
	.force_valid_4(force_valid_1_4_bottom_4),
	.force_valid_5(1'b0),

	.Arbitration_Result(Arbitration_1_4_bottom)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_2_1_mid
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(ref_force_valid[4]),
	.force_valid_1(force_valid_2_1_mid_1),
	.force_valid_2(force_valid_2_1_mid_2),
	.force_valid_3(force_valid_2_1_mid_3),
	.force_valid_4(force_valid_2_1_mid_4),
	.force_valid_5(force_valid_2_1_mid_5),

	.Arbitration_Result(Arbitration_2_1_mid)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_2_1_top
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_2_1_top_1),
	.force_valid_2(force_valid_2_1_top_2),
	.force_valid_3(force_valid_2_1_top_3),
	.force_valid_4(force_valid_2_1_top_4),
	.force_valid_5(force_valid_2_1_top_5),

	.Arbitration_Result(Arbitration_2_1_top)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_2_1_bottom
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_2_1_bottom_1),
	.force_valid_2(force_valid_2_1_bottom_2),
	.force_valid_3(force_valid_2_1_bottom_3),
	.force_valid_4(force_valid_2_1_bottom_4),
	.force_valid_5(1'b0),

	.Arbitration_Result(Arbitration_2_1_bottom)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_2_2_mid
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(ref_force_valid[5]),
	.force_valid_1(force_valid_2_2_mid_1),
	.force_valid_2(force_valid_2_2_mid_2),
	.force_valid_3(force_valid_2_2_mid_3),
	.force_valid_4(force_valid_2_2_mid_4),
	.force_valid_5(force_valid_2_2_mid_5),

	.Arbitration_Result(Arbitration_2_2_mid)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_2_2_top
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_2_2_top_1),
	.force_valid_2(force_valid_2_2_top_2),
	.force_valid_3(force_valid_2_2_top_3),
	.force_valid_4(force_valid_2_2_top_4),
	.force_valid_5(force_valid_2_2_top_5),

	.Arbitration_Result(Arbitration_2_2_top)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_2_2_bottom
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_2_2_bottom_1),
	.force_valid_2(force_valid_2_2_bottom_2),
	.force_valid_3(force_valid_2_2_bottom_3),
	.force_valid_4(force_valid_2_2_bottom_4),
	.force_valid_5(1'b0),

	.Arbitration_Result(Arbitration_2_2_bottom)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_2_3_mid
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(ref_force_valid[6]),
	.force_valid_1(force_valid_2_3_mid_1),
	.force_valid_2(force_valid_2_3_mid_2),
	.force_valid_3(force_valid_2_3_mid_3),
	.force_valid_4(force_valid_2_3_mid_4),
	.force_valid_5(force_valid_2_3_mid_5),

	.Arbitration_Result(Arbitration_2_3_mid)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_2_3_top
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_2_3_top_1),
	.force_valid_2(force_valid_2_3_top_2),
	.force_valid_3(force_valid_2_3_top_3),
	.force_valid_4(force_valid_2_3_top_4),
	.force_valid_5(force_valid_2_3_top_5),

	.Arbitration_Result(Arbitration_2_3_top)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_2_3_bottom
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_2_3_bottom_1),
	.force_valid_2(force_valid_2_3_bottom_2),
	.force_valid_3(force_valid_2_3_bottom_3),
	.force_valid_4(force_valid_2_3_bottom_4),
	.force_valid_5(1'b0),

	.Arbitration_Result(Arbitration_2_3_bottom)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_2_4_mid
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(ref_force_valid[7]),
	.force_valid_1(force_valid_2_4_mid_1),
	.force_valid_2(force_valid_2_4_mid_2),
	.force_valid_3(force_valid_2_4_mid_3),
	.force_valid_4(force_valid_2_4_mid_4),
	.force_valid_5(force_valid_2_4_mid_5),

	.Arbitration_Result(Arbitration_2_4_mid)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_2_4_top
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_2_4_top_1),
	.force_valid_2(force_valid_2_4_top_2),
	.force_valid_3(force_valid_2_4_top_3),
	.force_valid_4(force_valid_2_4_top_4),
	.force_valid_5(force_valid_2_4_top_5),

	.Arbitration_Result(Arbitration_2_4_top)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_2_4_bottom
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_2_4_bottom_1),
	.force_valid_2(force_valid_2_4_bottom_2),
	.force_valid_3(force_valid_2_4_bottom_3),
	.force_valid_4(force_valid_2_4_bottom_4),
	.force_valid_5(1'b0),

	.Arbitration_Result(Arbitration_2_4_bottom)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_3_1_mid
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(ref_force_valid[8]),
	.force_valid_1(force_valid_3_1_mid_1),
	.force_valid_2(force_valid_3_1_mid_2),
	.force_valid_3(force_valid_3_1_mid_3),
	.force_valid_4(force_valid_3_1_mid_4),
	.force_valid_5(force_valid_3_1_mid_5),

	.Arbitration_Result(Arbitration_3_1_mid)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_3_1_top
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_3_1_top_1),
	.force_valid_2(force_valid_3_1_top_2),
	.force_valid_3(force_valid_3_1_top_3),
	.force_valid_4(force_valid_3_1_top_4),
	.force_valid_5(force_valid_3_1_top_5),

	.Arbitration_Result(Arbitration_3_1_top)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_3_1_bottom
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_3_1_bottom_1),
	.force_valid_2(force_valid_3_1_bottom_2),
	.force_valid_3(force_valid_3_1_bottom_3),
	.force_valid_4(force_valid_3_1_bottom_4),
	.force_valid_5(1'b0),

	.Arbitration_Result(Arbitration_3_1_bottom)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_3_2_mid
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(ref_force_valid[9]),
	.force_valid_1(force_valid_3_2_mid_1),
	.force_valid_2(force_valid_3_2_mid_2),
	.force_valid_3(force_valid_3_2_mid_3),
	.force_valid_4(force_valid_3_2_mid_4),
	.force_valid_5(force_valid_3_2_mid_5),

	.Arbitration_Result(Arbitration_3_2_mid)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_3_2_top
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_3_2_top_1),
	.force_valid_2(force_valid_3_2_top_2),
	.force_valid_3(force_valid_3_2_top_3),
	.force_valid_4(force_valid_3_2_top_4),
	.force_valid_5(force_valid_3_2_top_5),

	.Arbitration_Result(Arbitration_3_2_top)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_3_2_bottom
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_3_2_bottom_1),
	.force_valid_2(force_valid_3_2_bottom_2),
	.force_valid_3(force_valid_3_2_bottom_3),
	.force_valid_4(force_valid_3_2_bottom_4),
	.force_valid_5(1'b0),

	.Arbitration_Result(Arbitration_3_2_bottom)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_3_3_mid
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(ref_force_valid[10]),
	.force_valid_1(force_valid_3_3_mid_1),
	.force_valid_2(force_valid_3_3_mid_2),
	.force_valid_3(force_valid_3_3_mid_3),
	.force_valid_4(force_valid_3_3_mid_4),
	.force_valid_5(force_valid_3_3_mid_5),

	.Arbitration_Result(Arbitration_3_3_mid)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_3_3_top
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_3_3_top_1),
	.force_valid_2(force_valid_3_3_top_2),
	.force_valid_3(force_valid_3_3_top_3),
	.force_valid_4(force_valid_3_3_top_4),
	.force_valid_5(force_valid_3_3_top_5),

	.Arbitration_Result(Arbitration_3_3_top)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_3_3_bottom
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_3_3_bottom_1),
	.force_valid_2(force_valid_3_3_bottom_2),
	.force_valid_3(force_valid_3_3_bottom_3),
	.force_valid_4(force_valid_3_3_bottom_4),
	.force_valid_5(1'b0),

	.Arbitration_Result(Arbitration_3_3_bottom)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_3_4_mid
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(ref_force_valid[11]),
	.force_valid_1(force_valid_3_4_mid_1),
	.force_valid_2(force_valid_3_4_mid_2),
	.force_valid_3(force_valid_3_4_mid_3),
	.force_valid_4(force_valid_3_4_mid_4),
	.force_valid_5(force_valid_3_4_mid_5),

	.Arbitration_Result(Arbitration_3_4_mid)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_3_4_top
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_3_4_top_1),
	.force_valid_2(force_valid_3_4_top_2),
	.force_valid_3(force_valid_3_4_top_3),
	.force_valid_4(force_valid_3_4_top_4),
	.force_valid_5(force_valid_3_4_top_5),

	.Arbitration_Result(Arbitration_3_4_top)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_3_4_bottom
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_3_4_bottom_1),
	.force_valid_2(force_valid_3_4_bottom_2),
	.force_valid_3(force_valid_3_4_bottom_3),
	.force_valid_4(force_valid_3_4_bottom_4),
	.force_valid_5(1'b0),

	.Arbitration_Result(Arbitration_3_4_bottom)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_4_1_mid
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(ref_force_valid[12]),
	.force_valid_1(force_valid_4_1_mid_1),
	.force_valid_2(force_valid_4_1_mid_2),
	.force_valid_3(force_valid_4_1_mid_3),
	.force_valid_4(force_valid_4_1_mid_4),
	.force_valid_5(force_valid_4_1_mid_5),

	.Arbitration_Result(Arbitration_4_1_mid)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_4_1_top
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_4_1_top_1),
	.force_valid_2(force_valid_4_1_top_2),
	.force_valid_3(force_valid_4_1_top_3),
	.force_valid_4(force_valid_4_1_top_4),
	.force_valid_5(force_valid_4_1_top_5),

	.Arbitration_Result(Arbitration_4_1_top)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_4_1_bottom
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_4_1_bottom_1),
	.force_valid_2(force_valid_4_1_bottom_2),
	.force_valid_3(force_valid_4_1_bottom_3),
	.force_valid_4(force_valid_4_1_bottom_4),
	.force_valid_5(1'b0),

	.Arbitration_Result(Arbitration_4_1_bottom)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_4_2_mid
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(ref_force_valid[13]),
	.force_valid_1(force_valid_4_2_mid_1),
	.force_valid_2(force_valid_4_2_mid_2),
	.force_valid_3(force_valid_4_2_mid_3),
	.force_valid_4(force_valid_4_2_mid_4),
	.force_valid_5(force_valid_4_2_mid_5),

	.Arbitration_Result(Arbitration_4_2_mid)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_4_2_top
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_4_2_top_1),
	.force_valid_2(force_valid_4_2_top_2),
	.force_valid_3(force_valid_4_2_top_3),
	.force_valid_4(force_valid_4_2_top_4),
	.force_valid_5(force_valid_4_2_top_5),

	.Arbitration_Result(Arbitration_4_2_top)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_4_2_bottom
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_4_2_bottom_1),
	.force_valid_2(force_valid_4_2_bottom_2),
	.force_valid_3(force_valid_4_2_bottom_3),
	.force_valid_4(force_valid_4_2_bottom_4),
	.force_valid_5(1'b0),

	.Arbitration_Result(Arbitration_4_2_bottom)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_4_3_mid
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(ref_force_valid[14]),
	.force_valid_1(force_valid_4_3_mid_1),
	.force_valid_2(force_valid_4_3_mid_2),
	.force_valid_3(force_valid_4_3_mid_3),
	.force_valid_4(force_valid_4_3_mid_4),
	.force_valid_5(force_valid_4_3_mid_5),

	.Arbitration_Result(Arbitration_4_3_mid)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_4_3_top
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_4_3_top_1),
	.force_valid_2(force_valid_4_3_top_2),
	.force_valid_3(force_valid_4_3_top_3),
	.force_valid_4(force_valid_4_3_top_4),
	.force_valid_5(force_valid_4_3_top_5),

	.Arbitration_Result(Arbitration_4_3_top)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_4_3_bottom
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_4_3_bottom_1),
	.force_valid_2(force_valid_4_3_bottom_2),
	.force_valid_3(force_valid_4_3_bottom_3),
	.force_valid_4(force_valid_4_3_bottom_4),
	.force_valid_5(1'b0),

	.Arbitration_Result(Arbitration_4_3_bottom)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_4_4_mid
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(ref_force_valid[15]),
	.force_valid_1(force_valid_4_4_mid_1),
	.force_valid_2(force_valid_4_4_mid_2),
	.force_valid_3(force_valid_4_4_mid_3),
	.force_valid_4(force_valid_4_4_mid_4),
	.force_valid_5(force_valid_4_4_mid_5),

	.Arbitration_Result(Arbitration_4_4_mid)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_4_4_top
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_4_4_top_1),
	.force_valid_2(force_valid_4_4_top_2),
	.force_valid_3(force_valid_4_4_top_3),
	.force_valid_4(force_valid_4_4_top_4),
	.force_valid_5(force_valid_4_4_top_5),

	.Arbitration_Result(Arbitration_4_4_top)
);
Force_Writeback_Arbiter
#(
	.FORCE_WTADDR_ARBITER_SIZE(FORCE_WTADDR_ARBITER_SIZE),
	.FORCE_WTADDR_ARBITER_MSB(FORCE_WTADDR_ARBITER_MSB)
)
Force_Writeback_Arbiter_4_4_bottom
(
	.clk(clk),
	.rst(rst),
	.ref_force_valid(1'b0),
	.force_valid_1(force_valid_4_4_bottom_1),
	.force_valid_2(force_valid_4_4_bottom_2),
	.force_valid_3(force_valid_4_4_bottom_3),
	.force_valid_4(force_valid_4_4_bottom_4),
	.force_valid_5(1'b0),

	.Arbitration_Result(Arbitration_4_4_bottom)
);

endmodule