/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Module: Mux_Tree.v
//
// Function: 
//				
//
// Data Organization:
//				
//
// Used by:
//				N/A
//
// Dependency:
//				N/A
//
// Testbench:
//				_tb.v
//
// Timing:
//				TBD
//
// Created by: 
//				Tong Geng 03/26/2019
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module Mux_Tree
#(
	parameter DATA_WIDTH 		= 32*3,
	parameter NUM_INPUT_PORTS	= 128,
	parameter SEL_DIWTH 		= $clog2(NUM_INPUT_PORTS)				// log(NUM_INPUT_PORTS) / log(2)
)
(
	input clk,
	input rst,
	input [SEL_DIWTH-1:0] in_sel,
	input [NUM_INPUT_PORTS-1:0] in_valid,
	input [NUM_INPUT_PORTS*DATA_WIDTH-1:0] in_data,
	output reg [DATA_WIDTH-1:0] out_data,
	output reg out_valid
);

    wire [NUM_INPUT_PORTS*DATA_WIDTH-1:0] in_data_reorder;
    reg [NUM_INPUT_PORTS*DATA_WIDTH-1:0] in_data_shifted;
    assign in_data_reorder = {in_data[12287],in_data[12191],in_data[12095],in_data[11999],in_data[11903],in_data[11807],in_data[11711],in_data[11615],in_data[11519],in_data[11423],in_data[11327],in_data[11231],in_data[11135],in_data[11039],in_data[10943],in_data[10847],in_data[10751],in_data[10655],in_data[10559],in_data[10463],in_data[10367],in_data[10271],in_data[10175],in_data[10079],in_data[9983],in_data[9887],in_data[9791],in_data[9695],in_data[9599],in_data[9503],in_data[9407],in_data[9311],in_data[9215],in_data[9119],in_data[9023],in_data[8927],in_data[8831],in_data[8735],in_data[8639],in_data[8543],in_data[8447],in_data[8351],in_data[8255],in_data[8159],in_data[8063],in_data[7967],in_data[7871],in_data[7775],in_data[7679],in_data[7583],in_data[7487],in_data[7391],in_data[7295],in_data[7199],in_data[7103],in_data[7007],in_data[6911],in_data[6815],in_data[6719],in_data[6623],in_data[6527],in_data[6431],in_data[6335],in_data[6239],in_data[6143],in_data[6047],in_data[5951],in_data[5855],in_data[5759],in_data[5663],in_data[5567],in_data[5471],in_data[5375],in_data[5279],in_data[5183],in_data[5087],in_data[4991],in_data[4895],in_data[4799],in_data[4703],in_data[4607],in_data[4511],in_data[4415],in_data[4319],in_data[4223],in_data[4127],in_data[4031],in_data[3935],in_data[3839],in_data[3743],in_data[3647],in_data[3551],in_data[3455],in_data[3359],in_data[3263],in_data[3167],in_data[3071],in_data[2975],in_data[2879],in_data[2783],in_data[2687],in_data[2591],in_data[2495],in_data[2399],in_data[2303],in_data[2207],in_data[2111],in_data[2015],in_data[1919],in_data[1823],in_data[1727],in_data[1631],in_data[1535],in_data[1439],in_data[1343],in_data[1247],in_data[1151],in_data[1055],in_data[959],in_data[863],in_data[767],in_data[671],in_data[575],in_data[479],in_data[383],in_data[287],in_data[191],in_data[95],in_data[12286],in_data[12190],in_data[12094],in_data[11998],in_data[11902],in_data[11806],in_data[11710],in_data[11614],in_data[11518],in_data[11422],in_data[11326],in_data[11230],in_data[11134],in_data[11038],in_data[10942],in_data[10846],in_data[10750],in_data[10654],in_data[10558],in_data[10462],in_data[10366],in_data[10270],in_data[10174],in_data[10078],in_data[9982],in_data[9886],in_data[9790],in_data[9694],in_data[9598],in_data[9502],in_data[9406],in_data[9310],in_data[9214],in_data[9118],in_data[9022],in_data[8926],in_data[8830],in_data[8734],in_data[8638],in_data[8542],in_data[8446],in_data[8350],in_data[8254],in_data[8158],in_data[8062],in_data[7966],in_data[7870],in_data[7774],in_data[7678],in_data[7582],in_data[7486],in_data[7390],in_data[7294],in_data[7198],in_data[7102],in_data[7006],in_data[6910],in_data[6814],in_data[6718],in_data[6622],in_data[6526],in_data[6430],in_data[6334],in_data[6238],in_data[6142],in_data[6046],in_data[5950],in_data[5854],in_data[5758],in_data[5662],in_data[5566],in_data[5470],in_data[5374],in_data[5278],in_data[5182],in_data[5086],in_data[4990],in_data[4894],in_data[4798],in_data[4702],in_data[4606],in_data[4510],in_data[4414],in_data[4318],in_data[4222],in_data[4126],in_data[4030],in_data[3934],in_data[3838],in_data[3742],in_data[3646],in_data[3550],in_data[3454],in_data[3358],in_data[3262],in_data[3166],in_data[3070],in_data[2974],in_data[2878],in_data[2782],in_data[2686],in_data[2590],in_data[2494],in_data[2398],in_data[2302],in_data[2206],in_data[2110],in_data[2014],in_data[1918],in_data[1822],in_data[1726],in_data[1630],in_data[1534],in_data[1438],in_data[1342],in_data[1246],in_data[1150],in_data[1054],in_data[958],in_data[862],in_data[766],in_data[670],in_data[574],in_data[478],in_data[382],in_data[286],in_data[190],in_data[94],in_data[12285],in_data[12189],in_data[12093],in_data[11997],in_data[11901],in_data[11805],in_data[11709],in_data[11613],in_data[11517],in_data[11421],in_data[11325],in_data[11229],in_data[11133],in_data[11037],in_data[10941],in_data[10845],in_data[10749],in_data[10653],in_data[10557],in_data[10461],in_data[10365],in_data[10269],in_data[10173],in_data[10077],in_data[9981],in_data[9885],in_data[9789],in_data[9693],in_data[9597],in_data[9501],in_data[9405],in_data[9309],in_data[9213],in_data[9117],in_data[9021],in_data[8925],in_data[8829],in_data[8733],in_data[8637],in_data[8541],in_data[8445],in_data[8349],in_data[8253],in_data[8157],in_data[8061],in_data[7965],in_data[7869],in_data[7773],in_data[7677],in_data[7581],in_data[7485],in_data[7389],in_data[7293],in_data[7197],in_data[7101],in_data[7005],in_data[6909],in_data[6813],in_data[6717],in_data[6621],in_data[6525],in_data[6429],in_data[6333],in_data[6237],in_data[6141],in_data[6045],in_data[5949],in_data[5853],in_data[5757],in_data[5661],in_data[5565],in_data[5469],in_data[5373],in_data[5277],in_data[5181],in_data[5085],in_data[4989],in_data[4893],in_data[4797],in_data[4701],in_data[4605],in_data[4509],in_data[4413],in_data[4317],in_data[4221],in_data[4125],in_data[4029],in_data[3933],in_data[3837],in_data[3741],in_data[3645],in_data[3549],in_data[3453],in_data[3357],in_data[3261],in_data[3165],in_data[3069],in_data[2973],in_data[2877],in_data[2781],in_data[2685],in_data[2589],in_data[2493],in_data[2397],in_data[2301],in_data[2205],in_data[2109],in_data[2013],in_data[1917],in_data[1821],in_data[1725],in_data[1629],in_data[1533],in_data[1437],in_data[1341],in_data[1245],in_data[1149],in_data[1053],in_data[957],in_data[861],in_data[765],in_data[669],in_data[573],in_data[477],in_data[381],in_data[285],in_data[189],in_data[93],in_data[12284],in_data[12188],in_data[12092],in_data[11996],in_data[11900],in_data[11804],in_data[11708],in_data[11612],in_data[11516],in_data[11420],in_data[11324],in_data[11228],in_data[11132],in_data[11036],in_data[10940],in_data[10844],in_data[10748],in_data[10652],in_data[10556],in_data[10460],in_data[10364],in_data[10268],in_data[10172],in_data[10076],in_data[9980],in_data[9884],in_data[9788],in_data[9692],in_data[9596],in_data[9500],in_data[9404],in_data[9308],in_data[9212],in_data[9116],in_data[9020],in_data[8924],in_data[8828],in_data[8732],in_data[8636],in_data[8540],in_data[8444],in_data[8348],in_data[8252],in_data[8156],in_data[8060],in_data[7964],in_data[7868],in_data[7772],in_data[7676],in_data[7580],in_data[7484],in_data[7388],in_data[7292],in_data[7196],in_data[7100],in_data[7004],in_data[6908],in_data[6812],in_data[6716],in_data[6620],in_data[6524],in_data[6428],in_data[6332],in_data[6236],in_data[6140],in_data[6044],in_data[5948],in_data[5852],in_data[5756],in_data[5660],in_data[5564],in_data[5468],in_data[5372],in_data[5276],in_data[5180],in_data[5084],in_data[4988],in_data[4892],in_data[4796],in_data[4700],in_data[4604],in_data[4508],in_data[4412],in_data[4316],in_data[4220],in_data[4124],in_data[4028],in_data[3932],in_data[3836],in_data[3740],in_data[3644],in_data[3548],in_data[3452],in_data[3356],in_data[3260],in_data[3164],in_data[3068],in_data[2972],in_data[2876],in_data[2780],in_data[2684],in_data[2588],in_data[2492],in_data[2396],in_data[2300],in_data[2204],in_data[2108],in_data[2012],in_data[1916],in_data[1820],in_data[1724],in_data[1628],in_data[1532],in_data[1436],in_data[1340],in_data[1244],in_data[1148],in_data[1052],in_data[956],in_data[860],in_data[764],in_data[668],in_data[572],in_data[476],in_data[380],in_data[284],in_data[188],in_data[92],in_data[12283],in_data[12187],in_data[12091],in_data[11995],in_data[11899],in_data[11803],in_data[11707],in_data[11611],in_data[11515],in_data[11419],in_data[11323],in_data[11227],in_data[11131],in_data[11035],in_data[10939],in_data[10843],in_data[10747],in_data[10651],in_data[10555],in_data[10459],in_data[10363],in_data[10267],in_data[10171],in_data[10075],in_data[9979],in_data[9883],in_data[9787],in_data[9691],in_data[9595],in_data[9499],in_data[9403],in_data[9307],in_data[9211],in_data[9115],in_data[9019],in_data[8923],in_data[8827],in_data[8731],in_data[8635],in_data[8539],in_data[8443],in_data[8347],in_data[8251],in_data[8155],in_data[8059],in_data[7963],in_data[7867],in_data[7771],in_data[7675],in_data[7579],in_data[7483],in_data[7387],in_data[7291],in_data[7195],in_data[7099],in_data[7003],in_data[6907],in_data[6811],in_data[6715],in_data[6619],in_data[6523],in_data[6427],in_data[6331],in_data[6235],in_data[6139],in_data[6043],in_data[5947],in_data[5851],in_data[5755],in_data[5659],in_data[5563],in_data[5467],in_data[5371],in_data[5275],in_data[5179],in_data[5083],in_data[4987],in_data[4891],in_data[4795],in_data[4699],in_data[4603],in_data[4507],in_data[4411],in_data[4315],in_data[4219],in_data[4123],in_data[4027],in_data[3931],in_data[3835],in_data[3739],in_data[3643],in_data[3547],in_data[3451],in_data[3355],in_data[3259],in_data[3163],in_data[3067],in_data[2971],in_data[2875],in_data[2779],in_data[2683],in_data[2587],in_data[2491],in_data[2395],in_data[2299],in_data[2203],in_data[2107],in_data[2011],in_data[1915],in_data[1819],in_data[1723],in_data[1627],in_data[1531],in_data[1435],in_data[1339],in_data[1243],in_data[1147],in_data[1051],in_data[955],in_data[859],in_data[763],in_data[667],in_data[571],in_data[475],in_data[379],in_data[283],in_data[187],in_data[91],in_data[12282],in_data[12186],in_data[12090],in_data[11994],in_data[11898],in_data[11802],in_data[11706],in_data[11610],in_data[11514],in_data[11418],in_data[11322],in_data[11226],in_data[11130],in_data[11034],in_data[10938],in_data[10842],in_data[10746],in_data[10650],in_data[10554],in_data[10458],in_data[10362],in_data[10266],in_data[10170],in_data[10074],in_data[9978],in_data[9882],in_data[9786],in_data[9690],in_data[9594],in_data[9498],in_data[9402],in_data[9306],in_data[9210],in_data[9114],in_data[9018],in_data[8922],in_data[8826],in_data[8730],in_data[8634],in_data[8538],in_data[8442],in_data[8346],in_data[8250],in_data[8154],in_data[8058],in_data[7962],in_data[7866],in_data[7770],in_data[7674],in_data[7578],in_data[7482],in_data[7386],in_data[7290],in_data[7194],in_data[7098],in_data[7002],in_data[6906],in_data[6810],in_data[6714],in_data[6618],in_data[6522],in_data[6426],in_data[6330],in_data[6234],in_data[6138],in_data[6042],in_data[5946],in_data[5850],in_data[5754],in_data[5658],in_data[5562],in_data[5466],in_data[5370],in_data[5274],in_data[5178],in_data[5082],in_data[4986],in_data[4890],in_data[4794],in_data[4698],in_data[4602],in_data[4506],in_data[4410],in_data[4314],in_data[4218],in_data[4122],in_data[4026],in_data[3930],in_data[3834],in_data[3738],in_data[3642],in_data[3546],in_data[3450],in_data[3354],in_data[3258],in_data[3162],in_data[3066],in_data[2970],in_data[2874],in_data[2778],in_data[2682],in_data[2586],in_data[2490],in_data[2394],in_data[2298],in_data[2202],in_data[2106],in_data[2010],in_data[1914],in_data[1818],in_data[1722],in_data[1626],in_data[1530],in_data[1434],in_data[1338],in_data[1242],in_data[1146],in_data[1050],in_data[954],in_data[858],in_data[762],in_data[666],in_data[570],in_data[474],in_data[378],in_data[282],in_data[186],in_data[90],in_data[12281],in_data[12185],in_data[12089],in_data[11993],in_data[11897],in_data[11801],in_data[11705],in_data[11609],in_data[11513],in_data[11417],in_data[11321],in_data[11225],in_data[11129],in_data[11033],in_data[10937],in_data[10841],in_data[10745],in_data[10649],in_data[10553],in_data[10457],in_data[10361],in_data[10265],in_data[10169],in_data[10073],in_data[9977],in_data[9881],in_data[9785],in_data[9689],in_data[9593],in_data[9497],in_data[9401],in_data[9305],in_data[9209],in_data[9113],in_data[9017],in_data[8921],in_data[8825],in_data[8729],in_data[8633],in_data[8537],in_data[8441],in_data[8345],in_data[8249],in_data[8153],in_data[8057],in_data[7961],in_data[7865],in_data[7769],in_data[7673],in_data[7577],in_data[7481],in_data[7385],in_data[7289],in_data[7193],in_data[7097],in_data[7001],in_data[6905],in_data[6809],in_data[6713],in_data[6617],in_data[6521],in_data[6425],in_data[6329],in_data[6233],in_data[6137],in_data[6041],in_data[5945],in_data[5849],in_data[5753],in_data[5657],in_data[5561],in_data[5465],in_data[5369],in_data[5273],in_data[5177],in_data[5081],in_data[4985],in_data[4889],in_data[4793],in_data[4697],in_data[4601],in_data[4505],in_data[4409],in_data[4313],in_data[4217],in_data[4121],in_data[4025],in_data[3929],in_data[3833],in_data[3737],in_data[3641],in_data[3545],in_data[3449],in_data[3353],in_data[3257],in_data[3161],in_data[3065],in_data[2969],in_data[2873],in_data[2777],in_data[2681],in_data[2585],in_data[2489],in_data[2393],in_data[2297],in_data[2201],in_data[2105],in_data[2009],in_data[1913],in_data[1817],in_data[1721],in_data[1625],in_data[1529],in_data[1433],in_data[1337],in_data[1241],in_data[1145],in_data[1049],in_data[953],in_data[857],in_data[761],in_data[665],in_data[569],in_data[473],in_data[377],in_data[281],in_data[185],in_data[89],in_data[12280],in_data[12184],in_data[12088],in_data[11992],in_data[11896],in_data[11800],in_data[11704],in_data[11608],in_data[11512],in_data[11416],in_data[11320],in_data[11224],in_data[11128],in_data[11032],in_data[10936],in_data[10840],in_data[10744],in_data[10648],in_data[10552],in_data[10456],in_data[10360],in_data[10264],in_data[10168],in_data[10072],in_data[9976],in_data[9880],in_data[9784],in_data[9688],in_data[9592],in_data[9496],in_data[9400],in_data[9304],in_data[9208],in_data[9112],in_data[9016],in_data[8920],in_data[8824],in_data[8728],in_data[8632],in_data[8536],in_data[8440],in_data[8344],in_data[8248],in_data[8152],in_data[8056],in_data[7960],in_data[7864],in_data[7768],in_data[7672],in_data[7576],in_data[7480],in_data[7384],in_data[7288],in_data[7192],in_data[7096],in_data[7000],in_data[6904],in_data[6808],in_data[6712],in_data[6616],in_data[6520],in_data[6424],in_data[6328],in_data[6232],in_data[6136],in_data[6040],in_data[5944],in_data[5848],in_data[5752],in_data[5656],in_data[5560],in_data[5464],in_data[5368],in_data[5272],in_data[5176],in_data[5080],in_data[4984],in_data[4888],in_data[4792],in_data[4696],in_data[4600],in_data[4504],in_data[4408],in_data[4312],in_data[4216],in_data[4120],in_data[4024],in_data[3928],in_data[3832],in_data[3736],in_data[3640],in_data[3544],in_data[3448],in_data[3352],in_data[3256],in_data[3160],in_data[3064],in_data[2968],in_data[2872],in_data[2776],in_data[2680],in_data[2584],in_data[2488],in_data[2392],in_data[2296],in_data[2200],in_data[2104],in_data[2008],in_data[1912],in_data[1816],in_data[1720],in_data[1624],in_data[1528],in_data[1432],in_data[1336],in_data[1240],in_data[1144],in_data[1048],in_data[952],in_data[856],in_data[760],in_data[664],in_data[568],in_data[472],in_data[376],in_data[280],in_data[184],in_data[88],in_data[12279],in_data[12183],in_data[12087],in_data[11991],in_data[11895],in_data[11799],in_data[11703],in_data[11607],in_data[11511],in_data[11415],in_data[11319],in_data[11223],in_data[11127],in_data[11031],in_data[10935],in_data[10839],in_data[10743],in_data[10647],in_data[10551],in_data[10455],in_data[10359],in_data[10263],in_data[10167],in_data[10071],in_data[9975],in_data[9879],in_data[9783],in_data[9687],in_data[9591],in_data[9495],in_data[9399],in_data[9303],in_data[9207],in_data[9111],in_data[9015],in_data[8919],in_data[8823],in_data[8727],in_data[8631],in_data[8535],in_data[8439],in_data[8343],in_data[8247],in_data[8151],in_data[8055],in_data[7959],in_data[7863],in_data[7767],in_data[7671],in_data[7575],in_data[7479],in_data[7383],in_data[7287],in_data[7191],in_data[7095],in_data[6999],in_data[6903],in_data[6807],in_data[6711],in_data[6615],in_data[6519],in_data[6423],in_data[6327],in_data[6231],in_data[6135],in_data[6039],in_data[5943],in_data[5847],in_data[5751],in_data[5655],in_data[5559],in_data[5463],in_data[5367],in_data[5271],in_data[5175],in_data[5079],in_data[4983],in_data[4887],in_data[4791],in_data[4695],in_data[4599],in_data[4503],in_data[4407],in_data[4311],in_data[4215],in_data[4119],in_data[4023],in_data[3927],in_data[3831],in_data[3735],in_data[3639],in_data[3543],in_data[3447],in_data[3351],in_data[3255],in_data[3159],in_data[3063],in_data[2967],in_data[2871],in_data[2775],in_data[2679],in_data[2583],in_data[2487],in_data[2391],in_data[2295],in_data[2199],in_data[2103],in_data[2007],in_data[1911],in_data[1815],in_data[1719],in_data[1623],in_data[1527],in_data[1431],in_data[1335],in_data[1239],in_data[1143],in_data[1047],in_data[951],in_data[855],in_data[759],in_data[663],in_data[567],in_data[471],in_data[375],in_data[279],in_data[183],in_data[87],in_data[12278],in_data[12182],in_data[12086],in_data[11990],in_data[11894],in_data[11798],in_data[11702],in_data[11606],in_data[11510],in_data[11414],in_data[11318],in_data[11222],in_data[11126],in_data[11030],in_data[10934],in_data[10838],in_data[10742],in_data[10646],in_data[10550],in_data[10454],in_data[10358],in_data[10262],in_data[10166],in_data[10070],in_data[9974],in_data[9878],in_data[9782],in_data[9686],in_data[9590],in_data[9494],in_data[9398],in_data[9302],in_data[9206],in_data[9110],in_data[9014],in_data[8918],in_data[8822],in_data[8726],in_data[8630],in_data[8534],in_data[8438],in_data[8342],in_data[8246],in_data[8150],in_data[8054],in_data[7958],in_data[7862],in_data[7766],in_data[7670],in_data[7574],in_data[7478],in_data[7382],in_data[7286],in_data[7190],in_data[7094],in_data[6998],in_data[6902],in_data[6806],in_data[6710],in_data[6614],in_data[6518],in_data[6422],in_data[6326],in_data[6230],in_data[6134],in_data[6038],in_data[5942],in_data[5846],in_data[5750],in_data[5654],in_data[5558],in_data[5462],in_data[5366],in_data[5270],in_data[5174],in_data[5078],in_data[4982],in_data[4886],in_data[4790],in_data[4694],in_data[4598],in_data[4502],in_data[4406],in_data[4310],in_data[4214],in_data[4118],in_data[4022],in_data[3926],in_data[3830],in_data[3734],in_data[3638],in_data[3542],in_data[3446],in_data[3350],in_data[3254],in_data[3158],in_data[3062],in_data[2966],in_data[2870],in_data[2774],in_data[2678],in_data[2582],in_data[2486],in_data[2390],in_data[2294],in_data[2198],in_data[2102],in_data[2006],in_data[1910],in_data[1814],in_data[1718],in_data[1622],in_data[1526],in_data[1430],in_data[1334],in_data[1238],in_data[1142],in_data[1046],in_data[950],in_data[854],in_data[758],in_data[662],in_data[566],in_data[470],in_data[374],in_data[278],in_data[182],in_data[86],in_data[12277],in_data[12181],in_data[12085],in_data[11989],in_data[11893],in_data[11797],in_data[11701],in_data[11605],in_data[11509],in_data[11413],in_data[11317],in_data[11221],in_data[11125],in_data[11029],in_data[10933],in_data[10837],in_data[10741],in_data[10645],in_data[10549],in_data[10453],in_data[10357],in_data[10261],in_data[10165],in_data[10069],in_data[9973],in_data[9877],in_data[9781],in_data[9685],in_data[9589],in_data[9493],in_data[9397],in_data[9301],in_data[9205],in_data[9109],in_data[9013],in_data[8917],in_data[8821],in_data[8725],in_data[8629],in_data[8533],in_data[8437],in_data[8341],in_data[8245],in_data[8149],in_data[8053],in_data[7957],in_data[7861],in_data[7765],in_data[7669],in_data[7573],in_data[7477],in_data[7381],in_data[7285],in_data[7189],in_data[7093],in_data[6997],in_data[6901],in_data[6805],in_data[6709],in_data[6613],in_data[6517],in_data[6421],in_data[6325],in_data[6229],in_data[6133],in_data[6037],in_data[5941],in_data[5845],in_data[5749],in_data[5653],in_data[5557],in_data[5461],in_data[5365],in_data[5269],in_data[5173],in_data[5077],in_data[4981],in_data[4885],in_data[4789],in_data[4693],in_data[4597],in_data[4501],in_data[4405],in_data[4309],in_data[4213],in_data[4117],in_data[4021],in_data[3925],in_data[3829],in_data[3733],in_data[3637],in_data[3541],in_data[3445],in_data[3349],in_data[3253],in_data[3157],in_data[3061],in_data[2965],in_data[2869],in_data[2773],in_data[2677],in_data[2581],in_data[2485],in_data[2389],in_data[2293],in_data[2197],in_data[2101],in_data[2005],in_data[1909],in_data[1813],in_data[1717],in_data[1621],in_data[1525],in_data[1429],in_data[1333],in_data[1237],in_data[1141],in_data[1045],in_data[949],in_data[853],in_data[757],in_data[661],in_data[565],in_data[469],in_data[373],in_data[277],in_data[181],in_data[85],in_data[12276],in_data[12180],in_data[12084],in_data[11988],in_data[11892],in_data[11796],in_data[11700],in_data[11604],in_data[11508],in_data[11412],in_data[11316],in_data[11220],in_data[11124],in_data[11028],in_data[10932],in_data[10836],in_data[10740],in_data[10644],in_data[10548],in_data[10452],in_data[10356],in_data[10260],in_data[10164],in_data[10068],in_data[9972],in_data[9876],in_data[9780],in_data[9684],in_data[9588],in_data[9492],in_data[9396],in_data[9300],in_data[9204],in_data[9108],in_data[9012],in_data[8916],in_data[8820],in_data[8724],in_data[8628],in_data[8532],in_data[8436],in_data[8340],in_data[8244],in_data[8148],in_data[8052],in_data[7956],in_data[7860],in_data[7764],in_data[7668],in_data[7572],in_data[7476],in_data[7380],in_data[7284],in_data[7188],in_data[7092],in_data[6996],in_data[6900],in_data[6804],in_data[6708],in_data[6612],in_data[6516],in_data[6420],in_data[6324],in_data[6228],in_data[6132],in_data[6036],in_data[5940],in_data[5844],in_data[5748],in_data[5652],in_data[5556],in_data[5460],in_data[5364],in_data[5268],in_data[5172],in_data[5076],in_data[4980],in_data[4884],in_data[4788],in_data[4692],in_data[4596],in_data[4500],in_data[4404],in_data[4308],in_data[4212],in_data[4116],in_data[4020],in_data[3924],in_data[3828],in_data[3732],in_data[3636],in_data[3540],in_data[3444],in_data[3348],in_data[3252],in_data[3156],in_data[3060],in_data[2964],in_data[2868],in_data[2772],in_data[2676],in_data[2580],in_data[2484],in_data[2388],in_data[2292],in_data[2196],in_data[2100],in_data[2004],in_data[1908],in_data[1812],in_data[1716],in_data[1620],in_data[1524],in_data[1428],in_data[1332],in_data[1236],in_data[1140],in_data[1044],in_data[948],in_data[852],in_data[756],in_data[660],in_data[564],in_data[468],in_data[372],in_data[276],in_data[180],in_data[84],in_data[12275],in_data[12179],in_data[12083],in_data[11987],in_data[11891],in_data[11795],in_data[11699],in_data[11603],in_data[11507],in_data[11411],in_data[11315],in_data[11219],in_data[11123],in_data[11027],in_data[10931],in_data[10835],in_data[10739],in_data[10643],in_data[10547],in_data[10451],in_data[10355],in_data[10259],in_data[10163],in_data[10067],in_data[9971],in_data[9875],in_data[9779],in_data[9683],in_data[9587],in_data[9491],in_data[9395],in_data[9299],in_data[9203],in_data[9107],in_data[9011],in_data[8915],in_data[8819],in_data[8723],in_data[8627],in_data[8531],in_data[8435],in_data[8339],in_data[8243],in_data[8147],in_data[8051],in_data[7955],in_data[7859],in_data[7763],in_data[7667],in_data[7571],in_data[7475],in_data[7379],in_data[7283],in_data[7187],in_data[7091],in_data[6995],in_data[6899],in_data[6803],in_data[6707],in_data[6611],in_data[6515],in_data[6419],in_data[6323],in_data[6227],in_data[6131],in_data[6035],in_data[5939],in_data[5843],in_data[5747],in_data[5651],in_data[5555],in_data[5459],in_data[5363],in_data[5267],in_data[5171],in_data[5075],in_data[4979],in_data[4883],in_data[4787],in_data[4691],in_data[4595],in_data[4499],in_data[4403],in_data[4307],in_data[4211],in_data[4115],in_data[4019],in_data[3923],in_data[3827],in_data[3731],in_data[3635],in_data[3539],in_data[3443],in_data[3347],in_data[3251],in_data[3155],in_data[3059],in_data[2963],in_data[2867],in_data[2771],in_data[2675],in_data[2579],in_data[2483],in_data[2387],in_data[2291],in_data[2195],in_data[2099],in_data[2003],in_data[1907],in_data[1811],in_data[1715],in_data[1619],in_data[1523],in_data[1427],in_data[1331],in_data[1235],in_data[1139],in_data[1043],in_data[947],in_data[851],in_data[755],in_data[659],in_data[563],in_data[467],in_data[371],in_data[275],in_data[179],in_data[83],in_data[12274],in_data[12178],in_data[12082],in_data[11986],in_data[11890],in_data[11794],in_data[11698],in_data[11602],in_data[11506],in_data[11410],in_data[11314],in_data[11218],in_data[11122],in_data[11026],in_data[10930],in_data[10834],in_data[10738],in_data[10642],in_data[10546],in_data[10450],in_data[10354],in_data[10258],in_data[10162],in_data[10066],in_data[9970],in_data[9874],in_data[9778],in_data[9682],in_data[9586],in_data[9490],in_data[9394],in_data[9298],in_data[9202],in_data[9106],in_data[9010],in_data[8914],in_data[8818],in_data[8722],in_data[8626],in_data[8530],in_data[8434],in_data[8338],in_data[8242],in_data[8146],in_data[8050],in_data[7954],in_data[7858],in_data[7762],in_data[7666],in_data[7570],in_data[7474],in_data[7378],in_data[7282],in_data[7186],in_data[7090],in_data[6994],in_data[6898],in_data[6802],in_data[6706],in_data[6610],in_data[6514],in_data[6418],in_data[6322],in_data[6226],in_data[6130],in_data[6034],in_data[5938],in_data[5842],in_data[5746],in_data[5650],in_data[5554],in_data[5458],in_data[5362],in_data[5266],in_data[5170],in_data[5074],in_data[4978],in_data[4882],in_data[4786],in_data[4690],in_data[4594],in_data[4498],in_data[4402],in_data[4306],in_data[4210],in_data[4114],in_data[4018],in_data[3922],in_data[3826],in_data[3730],in_data[3634],in_data[3538],in_data[3442],in_data[3346],in_data[3250],in_data[3154],in_data[3058],in_data[2962],in_data[2866],in_data[2770],in_data[2674],in_data[2578],in_data[2482],in_data[2386],in_data[2290],in_data[2194],in_data[2098],in_data[2002],in_data[1906],in_data[1810],in_data[1714],in_data[1618],in_data[1522],in_data[1426],in_data[1330],in_data[1234],in_data[1138],in_data[1042],in_data[946],in_data[850],in_data[754],in_data[658],in_data[562],in_data[466],in_data[370],in_data[274],in_data[178],in_data[82],in_data[12273],in_data[12177],in_data[12081],in_data[11985],in_data[11889],in_data[11793],in_data[11697],in_data[11601],in_data[11505],in_data[11409],in_data[11313],in_data[11217],in_data[11121],in_data[11025],in_data[10929],in_data[10833],in_data[10737],in_data[10641],in_data[10545],in_data[10449],in_data[10353],in_data[10257],in_data[10161],in_data[10065],in_data[9969],in_data[9873],in_data[9777],in_data[9681],in_data[9585],in_data[9489],in_data[9393],in_data[9297],in_data[9201],in_data[9105],in_data[9009],in_data[8913],in_data[8817],in_data[8721],in_data[8625],in_data[8529],in_data[8433],in_data[8337],in_data[8241],in_data[8145],in_data[8049],in_data[7953],in_data[7857],in_data[7761],in_data[7665],in_data[7569],in_data[7473],in_data[7377],in_data[7281],in_data[7185],in_data[7089],in_data[6993],in_data[6897],in_data[6801],in_data[6705],in_data[6609],in_data[6513],in_data[6417],in_data[6321],in_data[6225],in_data[6129],in_data[6033],in_data[5937],in_data[5841],in_data[5745],in_data[5649],in_data[5553],in_data[5457],in_data[5361],in_data[5265],in_data[5169],in_data[5073],in_data[4977],in_data[4881],in_data[4785],in_data[4689],in_data[4593],in_data[4497],in_data[4401],in_data[4305],in_data[4209],in_data[4113],in_data[4017],in_data[3921],in_data[3825],in_data[3729],in_data[3633],in_data[3537],in_data[3441],in_data[3345],in_data[3249],in_data[3153],in_data[3057],in_data[2961],in_data[2865],in_data[2769],in_data[2673],in_data[2577],in_data[2481],in_data[2385],in_data[2289],in_data[2193],in_data[2097],in_data[2001],in_data[1905],in_data[1809],in_data[1713],in_data[1617],in_data[1521],in_data[1425],in_data[1329],in_data[1233],in_data[1137],in_data[1041],in_data[945],in_data[849],in_data[753],in_data[657],in_data[561],in_data[465],in_data[369],in_data[273],in_data[177],in_data[81],in_data[12272],in_data[12176],in_data[12080],in_data[11984],in_data[11888],in_data[11792],in_data[11696],in_data[11600],in_data[11504],in_data[11408],in_data[11312],in_data[11216],in_data[11120],in_data[11024],in_data[10928],in_data[10832],in_data[10736],in_data[10640],in_data[10544],in_data[10448],in_data[10352],in_data[10256],in_data[10160],in_data[10064],in_data[9968],in_data[9872],in_data[9776],in_data[9680],in_data[9584],in_data[9488],in_data[9392],in_data[9296],in_data[9200],in_data[9104],in_data[9008],in_data[8912],in_data[8816],in_data[8720],in_data[8624],in_data[8528],in_data[8432],in_data[8336],in_data[8240],in_data[8144],in_data[8048],in_data[7952],in_data[7856],in_data[7760],in_data[7664],in_data[7568],in_data[7472],in_data[7376],in_data[7280],in_data[7184],in_data[7088],in_data[6992],in_data[6896],in_data[6800],in_data[6704],in_data[6608],in_data[6512],in_data[6416],in_data[6320],in_data[6224],in_data[6128],in_data[6032],in_data[5936],in_data[5840],in_data[5744],in_data[5648],in_data[5552],in_data[5456],in_data[5360],in_data[5264],in_data[5168],in_data[5072],in_data[4976],in_data[4880],in_data[4784],in_data[4688],in_data[4592],in_data[4496],in_data[4400],in_data[4304],in_data[4208],in_data[4112],in_data[4016],in_data[3920],in_data[3824],in_data[3728],in_data[3632],in_data[3536],in_data[3440],in_data[3344],in_data[3248],in_data[3152],in_data[3056],in_data[2960],in_data[2864],in_data[2768],in_data[2672],in_data[2576],in_data[2480],in_data[2384],in_data[2288],in_data[2192],in_data[2096],in_data[2000],in_data[1904],in_data[1808],in_data[1712],in_data[1616],in_data[1520],in_data[1424],in_data[1328],in_data[1232],in_data[1136],in_data[1040],in_data[944],in_data[848],in_data[752],in_data[656],in_data[560],in_data[464],in_data[368],in_data[272],in_data[176],in_data[80],in_data[12271],in_data[12175],in_data[12079],in_data[11983],in_data[11887],in_data[11791],in_data[11695],in_data[11599],in_data[11503],in_data[11407],in_data[11311],in_data[11215],in_data[11119],in_data[11023],in_data[10927],in_data[10831],in_data[10735],in_data[10639],in_data[10543],in_data[10447],in_data[10351],in_data[10255],in_data[10159],in_data[10063],in_data[9967],in_data[9871],in_data[9775],in_data[9679],in_data[9583],in_data[9487],in_data[9391],in_data[9295],in_data[9199],in_data[9103],in_data[9007],in_data[8911],in_data[8815],in_data[8719],in_data[8623],in_data[8527],in_data[8431],in_data[8335],in_data[8239],in_data[8143],in_data[8047],in_data[7951],in_data[7855],in_data[7759],in_data[7663],in_data[7567],in_data[7471],in_data[7375],in_data[7279],in_data[7183],in_data[7087],in_data[6991],in_data[6895],in_data[6799],in_data[6703],in_data[6607],in_data[6511],in_data[6415],in_data[6319],in_data[6223],in_data[6127],in_data[6031],in_data[5935],in_data[5839],in_data[5743],in_data[5647],in_data[5551],in_data[5455],in_data[5359],in_data[5263],in_data[5167],in_data[5071],in_data[4975],in_data[4879],in_data[4783],in_data[4687],in_data[4591],in_data[4495],in_data[4399],in_data[4303],in_data[4207],in_data[4111],in_data[4015],in_data[3919],in_data[3823],in_data[3727],in_data[3631],in_data[3535],in_data[3439],in_data[3343],in_data[3247],in_data[3151],in_data[3055],in_data[2959],in_data[2863],in_data[2767],in_data[2671],in_data[2575],in_data[2479],in_data[2383],in_data[2287],in_data[2191],in_data[2095],in_data[1999],in_data[1903],in_data[1807],in_data[1711],in_data[1615],in_data[1519],in_data[1423],in_data[1327],in_data[1231],in_data[1135],in_data[1039],in_data[943],in_data[847],in_data[751],in_data[655],in_data[559],in_data[463],in_data[367],in_data[271],in_data[175],in_data[79],in_data[12270],in_data[12174],in_data[12078],in_data[11982],in_data[11886],in_data[11790],in_data[11694],in_data[11598],in_data[11502],in_data[11406],in_data[11310],in_data[11214],in_data[11118],in_data[11022],in_data[10926],in_data[10830],in_data[10734],in_data[10638],in_data[10542],in_data[10446],in_data[10350],in_data[10254],in_data[10158],in_data[10062],in_data[9966],in_data[9870],in_data[9774],in_data[9678],in_data[9582],in_data[9486],in_data[9390],in_data[9294],in_data[9198],in_data[9102],in_data[9006],in_data[8910],in_data[8814],in_data[8718],in_data[8622],in_data[8526],in_data[8430],in_data[8334],in_data[8238],in_data[8142],in_data[8046],in_data[7950],in_data[7854],in_data[7758],in_data[7662],in_data[7566],in_data[7470],in_data[7374],in_data[7278],in_data[7182],in_data[7086],in_data[6990],in_data[6894],in_data[6798],in_data[6702],in_data[6606],in_data[6510],in_data[6414],in_data[6318],in_data[6222],in_data[6126],in_data[6030],in_data[5934],in_data[5838],in_data[5742],in_data[5646],in_data[5550],in_data[5454],in_data[5358],in_data[5262],in_data[5166],in_data[5070],in_data[4974],in_data[4878],in_data[4782],in_data[4686],in_data[4590],in_data[4494],in_data[4398],in_data[4302],in_data[4206],in_data[4110],in_data[4014],in_data[3918],in_data[3822],in_data[3726],in_data[3630],in_data[3534],in_data[3438],in_data[3342],in_data[3246],in_data[3150],in_data[3054],in_data[2958],in_data[2862],in_data[2766],in_data[2670],in_data[2574],in_data[2478],in_data[2382],in_data[2286],in_data[2190],in_data[2094],in_data[1998],in_data[1902],in_data[1806],in_data[1710],in_data[1614],in_data[1518],in_data[1422],in_data[1326],in_data[1230],in_data[1134],in_data[1038],in_data[942],in_data[846],in_data[750],in_data[654],in_data[558],in_data[462],in_data[366],in_data[270],in_data[174],in_data[78],in_data[12269],in_data[12173],in_data[12077],in_data[11981],in_data[11885],in_data[11789],in_data[11693],in_data[11597],in_data[11501],in_data[11405],in_data[11309],in_data[11213],in_data[11117],in_data[11021],in_data[10925],in_data[10829],in_data[10733],in_data[10637],in_data[10541],in_data[10445],in_data[10349],in_data[10253],in_data[10157],in_data[10061],in_data[9965],in_data[9869],in_data[9773],in_data[9677],in_data[9581],in_data[9485],in_data[9389],in_data[9293],in_data[9197],in_data[9101],in_data[9005],in_data[8909],in_data[8813],in_data[8717],in_data[8621],in_data[8525],in_data[8429],in_data[8333],in_data[8237],in_data[8141],in_data[8045],in_data[7949],in_data[7853],in_data[7757],in_data[7661],in_data[7565],in_data[7469],in_data[7373],in_data[7277],in_data[7181],in_data[7085],in_data[6989],in_data[6893],in_data[6797],in_data[6701],in_data[6605],in_data[6509],in_data[6413],in_data[6317],in_data[6221],in_data[6125],in_data[6029],in_data[5933],in_data[5837],in_data[5741],in_data[5645],in_data[5549],in_data[5453],in_data[5357],in_data[5261],in_data[5165],in_data[5069],in_data[4973],in_data[4877],in_data[4781],in_data[4685],in_data[4589],in_data[4493],in_data[4397],in_data[4301],in_data[4205],in_data[4109],in_data[4013],in_data[3917],in_data[3821],in_data[3725],in_data[3629],in_data[3533],in_data[3437],in_data[3341],in_data[3245],in_data[3149],in_data[3053],in_data[2957],in_data[2861],in_data[2765],in_data[2669],in_data[2573],in_data[2477],in_data[2381],in_data[2285],in_data[2189],in_data[2093],in_data[1997],in_data[1901],in_data[1805],in_data[1709],in_data[1613],in_data[1517],in_data[1421],in_data[1325],in_data[1229],in_data[1133],in_data[1037],in_data[941],in_data[845],in_data[749],in_data[653],in_data[557],in_data[461],in_data[365],in_data[269],in_data[173],in_data[77],in_data[12268],in_data[12172],in_data[12076],in_data[11980],in_data[11884],in_data[11788],in_data[11692],in_data[11596],in_data[11500],in_data[11404],in_data[11308],in_data[11212],in_data[11116],in_data[11020],in_data[10924],in_data[10828],in_data[10732],in_data[10636],in_data[10540],in_data[10444],in_data[10348],in_data[10252],in_data[10156],in_data[10060],in_data[9964],in_data[9868],in_data[9772],in_data[9676],in_data[9580],in_data[9484],in_data[9388],in_data[9292],in_data[9196],in_data[9100],in_data[9004],in_data[8908],in_data[8812],in_data[8716],in_data[8620],in_data[8524],in_data[8428],in_data[8332],in_data[8236],in_data[8140],in_data[8044],in_data[7948],in_data[7852],in_data[7756],in_data[7660],in_data[7564],in_data[7468],in_data[7372],in_data[7276],in_data[7180],in_data[7084],in_data[6988],in_data[6892],in_data[6796],in_data[6700],in_data[6604],in_data[6508],in_data[6412],in_data[6316],in_data[6220],in_data[6124],in_data[6028],in_data[5932],in_data[5836],in_data[5740],in_data[5644],in_data[5548],in_data[5452],in_data[5356],in_data[5260],in_data[5164],in_data[5068],in_data[4972],in_data[4876],in_data[4780],in_data[4684],in_data[4588],in_data[4492],in_data[4396],in_data[4300],in_data[4204],in_data[4108],in_data[4012],in_data[3916],in_data[3820],in_data[3724],in_data[3628],in_data[3532],in_data[3436],in_data[3340],in_data[3244],in_data[3148],in_data[3052],in_data[2956],in_data[2860],in_data[2764],in_data[2668],in_data[2572],in_data[2476],in_data[2380],in_data[2284],in_data[2188],in_data[2092],in_data[1996],in_data[1900],in_data[1804],in_data[1708],in_data[1612],in_data[1516],in_data[1420],in_data[1324],in_data[1228],in_data[1132],in_data[1036],in_data[940],in_data[844],in_data[748],in_data[652],in_data[556],in_data[460],in_data[364],in_data[268],in_data[172],in_data[76],in_data[12267],in_data[12171],in_data[12075],in_data[11979],in_data[11883],in_data[11787],in_data[11691],in_data[11595],in_data[11499],in_data[11403],in_data[11307],in_data[11211],in_data[11115],in_data[11019],in_data[10923],in_data[10827],in_data[10731],in_data[10635],in_data[10539],in_data[10443],in_data[10347],in_data[10251],in_data[10155],in_data[10059],in_data[9963],in_data[9867],in_data[9771],in_data[9675],in_data[9579],in_data[9483],in_data[9387],in_data[9291],in_data[9195],in_data[9099],in_data[9003],in_data[8907],in_data[8811],in_data[8715],in_data[8619],in_data[8523],in_data[8427],in_data[8331],in_data[8235],in_data[8139],in_data[8043],in_data[7947],in_data[7851],in_data[7755],in_data[7659],in_data[7563],in_data[7467],in_data[7371],in_data[7275],in_data[7179],in_data[7083],in_data[6987],in_data[6891],in_data[6795],in_data[6699],in_data[6603],in_data[6507],in_data[6411],in_data[6315],in_data[6219],in_data[6123],in_data[6027],in_data[5931],in_data[5835],in_data[5739],in_data[5643],in_data[5547],in_data[5451],in_data[5355],in_data[5259],in_data[5163],in_data[5067],in_data[4971],in_data[4875],in_data[4779],in_data[4683],in_data[4587],in_data[4491],in_data[4395],in_data[4299],in_data[4203],in_data[4107],in_data[4011],in_data[3915],in_data[3819],in_data[3723],in_data[3627],in_data[3531],in_data[3435],in_data[3339],in_data[3243],in_data[3147],in_data[3051],in_data[2955],in_data[2859],in_data[2763],in_data[2667],in_data[2571],in_data[2475],in_data[2379],in_data[2283],in_data[2187],in_data[2091],in_data[1995],in_data[1899],in_data[1803],in_data[1707],in_data[1611],in_data[1515],in_data[1419],in_data[1323],in_data[1227],in_data[1131],in_data[1035],in_data[939],in_data[843],in_data[747],in_data[651],in_data[555],in_data[459],in_data[363],in_data[267],in_data[171],in_data[75],in_data[12266],in_data[12170],in_data[12074],in_data[11978],in_data[11882],in_data[11786],in_data[11690],in_data[11594],in_data[11498],in_data[11402],in_data[11306],in_data[11210],in_data[11114],in_data[11018],in_data[10922],in_data[10826],in_data[10730],in_data[10634],in_data[10538],in_data[10442],in_data[10346],in_data[10250],in_data[10154],in_data[10058],in_data[9962],in_data[9866],in_data[9770],in_data[9674],in_data[9578],in_data[9482],in_data[9386],in_data[9290],in_data[9194],in_data[9098],in_data[9002],in_data[8906],in_data[8810],in_data[8714],in_data[8618],in_data[8522],in_data[8426],in_data[8330],in_data[8234],in_data[8138],in_data[8042],in_data[7946],in_data[7850],in_data[7754],in_data[7658],in_data[7562],in_data[7466],in_data[7370],in_data[7274],in_data[7178],in_data[7082],in_data[6986],in_data[6890],in_data[6794],in_data[6698],in_data[6602],in_data[6506],in_data[6410],in_data[6314],in_data[6218],in_data[6122],in_data[6026],in_data[5930],in_data[5834],in_data[5738],in_data[5642],in_data[5546],in_data[5450],in_data[5354],in_data[5258],in_data[5162],in_data[5066],in_data[4970],in_data[4874],in_data[4778],in_data[4682],in_data[4586],in_data[4490],in_data[4394],in_data[4298],in_data[4202],in_data[4106],in_data[4010],in_data[3914],in_data[3818],in_data[3722],in_data[3626],in_data[3530],in_data[3434],in_data[3338],in_data[3242],in_data[3146],in_data[3050],in_data[2954],in_data[2858],in_data[2762],in_data[2666],in_data[2570],in_data[2474],in_data[2378],in_data[2282],in_data[2186],in_data[2090],in_data[1994],in_data[1898],in_data[1802],in_data[1706],in_data[1610],in_data[1514],in_data[1418],in_data[1322],in_data[1226],in_data[1130],in_data[1034],in_data[938],in_data[842],in_data[746],in_data[650],in_data[554],in_data[458],in_data[362],in_data[266],in_data[170],in_data[74],in_data[12265],in_data[12169],in_data[12073],in_data[11977],in_data[11881],in_data[11785],in_data[11689],in_data[11593],in_data[11497],in_data[11401],in_data[11305],in_data[11209],in_data[11113],in_data[11017],in_data[10921],in_data[10825],in_data[10729],in_data[10633],in_data[10537],in_data[10441],in_data[10345],in_data[10249],in_data[10153],in_data[10057],in_data[9961],in_data[9865],in_data[9769],in_data[9673],in_data[9577],in_data[9481],in_data[9385],in_data[9289],in_data[9193],in_data[9097],in_data[9001],in_data[8905],in_data[8809],in_data[8713],in_data[8617],in_data[8521],in_data[8425],in_data[8329],in_data[8233],in_data[8137],in_data[8041],in_data[7945],in_data[7849],in_data[7753],in_data[7657],in_data[7561],in_data[7465],in_data[7369],in_data[7273],in_data[7177],in_data[7081],in_data[6985],in_data[6889],in_data[6793],in_data[6697],in_data[6601],in_data[6505],in_data[6409],in_data[6313],in_data[6217],in_data[6121],in_data[6025],in_data[5929],in_data[5833],in_data[5737],in_data[5641],in_data[5545],in_data[5449],in_data[5353],in_data[5257],in_data[5161],in_data[5065],in_data[4969],in_data[4873],in_data[4777],in_data[4681],in_data[4585],in_data[4489],in_data[4393],in_data[4297],in_data[4201],in_data[4105],in_data[4009],in_data[3913],in_data[3817],in_data[3721],in_data[3625],in_data[3529],in_data[3433],in_data[3337],in_data[3241],in_data[3145],in_data[3049],in_data[2953],in_data[2857],in_data[2761],in_data[2665],in_data[2569],in_data[2473],in_data[2377],in_data[2281],in_data[2185],in_data[2089],in_data[1993],in_data[1897],in_data[1801],in_data[1705],in_data[1609],in_data[1513],in_data[1417],in_data[1321],in_data[1225],in_data[1129],in_data[1033],in_data[937],in_data[841],in_data[745],in_data[649],in_data[553],in_data[457],in_data[361],in_data[265],in_data[169],in_data[73],in_data[12264],in_data[12168],in_data[12072],in_data[11976],in_data[11880],in_data[11784],in_data[11688],in_data[11592],in_data[11496],in_data[11400],in_data[11304],in_data[11208],in_data[11112],in_data[11016],in_data[10920],in_data[10824],in_data[10728],in_data[10632],in_data[10536],in_data[10440],in_data[10344],in_data[10248],in_data[10152],in_data[10056],in_data[9960],in_data[9864],in_data[9768],in_data[9672],in_data[9576],in_data[9480],in_data[9384],in_data[9288],in_data[9192],in_data[9096],in_data[9000],in_data[8904],in_data[8808],in_data[8712],in_data[8616],in_data[8520],in_data[8424],in_data[8328],in_data[8232],in_data[8136],in_data[8040],in_data[7944],in_data[7848],in_data[7752],in_data[7656],in_data[7560],in_data[7464],in_data[7368],in_data[7272],in_data[7176],in_data[7080],in_data[6984],in_data[6888],in_data[6792],in_data[6696],in_data[6600],in_data[6504],in_data[6408],in_data[6312],in_data[6216],in_data[6120],in_data[6024],in_data[5928],in_data[5832],in_data[5736],in_data[5640],in_data[5544],in_data[5448],in_data[5352],in_data[5256],in_data[5160],in_data[5064],in_data[4968],in_data[4872],in_data[4776],in_data[4680],in_data[4584],in_data[4488],in_data[4392],in_data[4296],in_data[4200],in_data[4104],in_data[4008],in_data[3912],in_data[3816],in_data[3720],in_data[3624],in_data[3528],in_data[3432],in_data[3336],in_data[3240],in_data[3144],in_data[3048],in_data[2952],in_data[2856],in_data[2760],in_data[2664],in_data[2568],in_data[2472],in_data[2376],in_data[2280],in_data[2184],in_data[2088],in_data[1992],in_data[1896],in_data[1800],in_data[1704],in_data[1608],in_data[1512],in_data[1416],in_data[1320],in_data[1224],in_data[1128],in_data[1032],in_data[936],in_data[840],in_data[744],in_data[648],in_data[552],in_data[456],in_data[360],in_data[264],in_data[168],in_data[72],in_data[12263],in_data[12167],in_data[12071],in_data[11975],in_data[11879],in_data[11783],in_data[11687],in_data[11591],in_data[11495],in_data[11399],in_data[11303],in_data[11207],in_data[11111],in_data[11015],in_data[10919],in_data[10823],in_data[10727],in_data[10631],in_data[10535],in_data[10439],in_data[10343],in_data[10247],in_data[10151],in_data[10055],in_data[9959],in_data[9863],in_data[9767],in_data[9671],in_data[9575],in_data[9479],in_data[9383],in_data[9287],in_data[9191],in_data[9095],in_data[8999],in_data[8903],in_data[8807],in_data[8711],in_data[8615],in_data[8519],in_data[8423],in_data[8327],in_data[8231],in_data[8135],in_data[8039],in_data[7943],in_data[7847],in_data[7751],in_data[7655],in_data[7559],in_data[7463],in_data[7367],in_data[7271],in_data[7175],in_data[7079],in_data[6983],in_data[6887],in_data[6791],in_data[6695],in_data[6599],in_data[6503],in_data[6407],in_data[6311],in_data[6215],in_data[6119],in_data[6023],in_data[5927],in_data[5831],in_data[5735],in_data[5639],in_data[5543],in_data[5447],in_data[5351],in_data[5255],in_data[5159],in_data[5063],in_data[4967],in_data[4871],in_data[4775],in_data[4679],in_data[4583],in_data[4487],in_data[4391],in_data[4295],in_data[4199],in_data[4103],in_data[4007],in_data[3911],in_data[3815],in_data[3719],in_data[3623],in_data[3527],in_data[3431],in_data[3335],in_data[3239],in_data[3143],in_data[3047],in_data[2951],in_data[2855],in_data[2759],in_data[2663],in_data[2567],in_data[2471],in_data[2375],in_data[2279],in_data[2183],in_data[2087],in_data[1991],in_data[1895],in_data[1799],in_data[1703],in_data[1607],in_data[1511],in_data[1415],in_data[1319],in_data[1223],in_data[1127],in_data[1031],in_data[935],in_data[839],in_data[743],in_data[647],in_data[551],in_data[455],in_data[359],in_data[263],in_data[167],in_data[71],in_data[12262],in_data[12166],in_data[12070],in_data[11974],in_data[11878],in_data[11782],in_data[11686],in_data[11590],in_data[11494],in_data[11398],in_data[11302],in_data[11206],in_data[11110],in_data[11014],in_data[10918],in_data[10822],in_data[10726],in_data[10630],in_data[10534],in_data[10438],in_data[10342],in_data[10246],in_data[10150],in_data[10054],in_data[9958],in_data[9862],in_data[9766],in_data[9670],in_data[9574],in_data[9478],in_data[9382],in_data[9286],in_data[9190],in_data[9094],in_data[8998],in_data[8902],in_data[8806],in_data[8710],in_data[8614],in_data[8518],in_data[8422],in_data[8326],in_data[8230],in_data[8134],in_data[8038],in_data[7942],in_data[7846],in_data[7750],in_data[7654],in_data[7558],in_data[7462],in_data[7366],in_data[7270],in_data[7174],in_data[7078],in_data[6982],in_data[6886],in_data[6790],in_data[6694],in_data[6598],in_data[6502],in_data[6406],in_data[6310],in_data[6214],in_data[6118],in_data[6022],in_data[5926],in_data[5830],in_data[5734],in_data[5638],in_data[5542],in_data[5446],in_data[5350],in_data[5254],in_data[5158],in_data[5062],in_data[4966],in_data[4870],in_data[4774],in_data[4678],in_data[4582],in_data[4486],in_data[4390],in_data[4294],in_data[4198],in_data[4102],in_data[4006],in_data[3910],in_data[3814],in_data[3718],in_data[3622],in_data[3526],in_data[3430],in_data[3334],in_data[3238],in_data[3142],in_data[3046],in_data[2950],in_data[2854],in_data[2758],in_data[2662],in_data[2566],in_data[2470],in_data[2374],in_data[2278],in_data[2182],in_data[2086],in_data[1990],in_data[1894],in_data[1798],in_data[1702],in_data[1606],in_data[1510],in_data[1414],in_data[1318],in_data[1222],in_data[1126],in_data[1030],in_data[934],in_data[838],in_data[742],in_data[646],in_data[550],in_data[454],in_data[358],in_data[262],in_data[166],in_data[70],in_data[12261],in_data[12165],in_data[12069],in_data[11973],in_data[11877],in_data[11781],in_data[11685],in_data[11589],in_data[11493],in_data[11397],in_data[11301],in_data[11205],in_data[11109],in_data[11013],in_data[10917],in_data[10821],in_data[10725],in_data[10629],in_data[10533],in_data[10437],in_data[10341],in_data[10245],in_data[10149],in_data[10053],in_data[9957],in_data[9861],in_data[9765],in_data[9669],in_data[9573],in_data[9477],in_data[9381],in_data[9285],in_data[9189],in_data[9093],in_data[8997],in_data[8901],in_data[8805],in_data[8709],in_data[8613],in_data[8517],in_data[8421],in_data[8325],in_data[8229],in_data[8133],in_data[8037],in_data[7941],in_data[7845],in_data[7749],in_data[7653],in_data[7557],in_data[7461],in_data[7365],in_data[7269],in_data[7173],in_data[7077],in_data[6981],in_data[6885],in_data[6789],in_data[6693],in_data[6597],in_data[6501],in_data[6405],in_data[6309],in_data[6213],in_data[6117],in_data[6021],in_data[5925],in_data[5829],in_data[5733],in_data[5637],in_data[5541],in_data[5445],in_data[5349],in_data[5253],in_data[5157],in_data[5061],in_data[4965],in_data[4869],in_data[4773],in_data[4677],in_data[4581],in_data[4485],in_data[4389],in_data[4293],in_data[4197],in_data[4101],in_data[4005],in_data[3909],in_data[3813],in_data[3717],in_data[3621],in_data[3525],in_data[3429],in_data[3333],in_data[3237],in_data[3141],in_data[3045],in_data[2949],in_data[2853],in_data[2757],in_data[2661],in_data[2565],in_data[2469],in_data[2373],in_data[2277],in_data[2181],in_data[2085],in_data[1989],in_data[1893],in_data[1797],in_data[1701],in_data[1605],in_data[1509],in_data[1413],in_data[1317],in_data[1221],in_data[1125],in_data[1029],in_data[933],in_data[837],in_data[741],in_data[645],in_data[549],in_data[453],in_data[357],in_data[261],in_data[165],in_data[69],in_data[12260],in_data[12164],in_data[12068],in_data[11972],in_data[11876],in_data[11780],in_data[11684],in_data[11588],in_data[11492],in_data[11396],in_data[11300],in_data[11204],in_data[11108],in_data[11012],in_data[10916],in_data[10820],in_data[10724],in_data[10628],in_data[10532],in_data[10436],in_data[10340],in_data[10244],in_data[10148],in_data[10052],in_data[9956],in_data[9860],in_data[9764],in_data[9668],in_data[9572],in_data[9476],in_data[9380],in_data[9284],in_data[9188],in_data[9092],in_data[8996],in_data[8900],in_data[8804],in_data[8708],in_data[8612],in_data[8516],in_data[8420],in_data[8324],in_data[8228],in_data[8132],in_data[8036],in_data[7940],in_data[7844],in_data[7748],in_data[7652],in_data[7556],in_data[7460],in_data[7364],in_data[7268],in_data[7172],in_data[7076],in_data[6980],in_data[6884],in_data[6788],in_data[6692],in_data[6596],in_data[6500],in_data[6404],in_data[6308],in_data[6212],in_data[6116],in_data[6020],in_data[5924],in_data[5828],in_data[5732],in_data[5636],in_data[5540],in_data[5444],in_data[5348],in_data[5252],in_data[5156],in_data[5060],in_data[4964],in_data[4868],in_data[4772],in_data[4676],in_data[4580],in_data[4484],in_data[4388],in_data[4292],in_data[4196],in_data[4100],in_data[4004],in_data[3908],in_data[3812],in_data[3716],in_data[3620],in_data[3524],in_data[3428],in_data[3332],in_data[3236],in_data[3140],in_data[3044],in_data[2948],in_data[2852],in_data[2756],in_data[2660],in_data[2564],in_data[2468],in_data[2372],in_data[2276],in_data[2180],in_data[2084],in_data[1988],in_data[1892],in_data[1796],in_data[1700],in_data[1604],in_data[1508],in_data[1412],in_data[1316],in_data[1220],in_data[1124],in_data[1028],in_data[932],in_data[836],in_data[740],in_data[644],in_data[548],in_data[452],in_data[356],in_data[260],in_data[164],in_data[68],in_data[12259],in_data[12163],in_data[12067],in_data[11971],in_data[11875],in_data[11779],in_data[11683],in_data[11587],in_data[11491],in_data[11395],in_data[11299],in_data[11203],in_data[11107],in_data[11011],in_data[10915],in_data[10819],in_data[10723],in_data[10627],in_data[10531],in_data[10435],in_data[10339],in_data[10243],in_data[10147],in_data[10051],in_data[9955],in_data[9859],in_data[9763],in_data[9667],in_data[9571],in_data[9475],in_data[9379],in_data[9283],in_data[9187],in_data[9091],in_data[8995],in_data[8899],in_data[8803],in_data[8707],in_data[8611],in_data[8515],in_data[8419],in_data[8323],in_data[8227],in_data[8131],in_data[8035],in_data[7939],in_data[7843],in_data[7747],in_data[7651],in_data[7555],in_data[7459],in_data[7363],in_data[7267],in_data[7171],in_data[7075],in_data[6979],in_data[6883],in_data[6787],in_data[6691],in_data[6595],in_data[6499],in_data[6403],in_data[6307],in_data[6211],in_data[6115],in_data[6019],in_data[5923],in_data[5827],in_data[5731],in_data[5635],in_data[5539],in_data[5443],in_data[5347],in_data[5251],in_data[5155],in_data[5059],in_data[4963],in_data[4867],in_data[4771],in_data[4675],in_data[4579],in_data[4483],in_data[4387],in_data[4291],in_data[4195],in_data[4099],in_data[4003],in_data[3907],in_data[3811],in_data[3715],in_data[3619],in_data[3523],in_data[3427],in_data[3331],in_data[3235],in_data[3139],in_data[3043],in_data[2947],in_data[2851],in_data[2755],in_data[2659],in_data[2563],in_data[2467],in_data[2371],in_data[2275],in_data[2179],in_data[2083],in_data[1987],in_data[1891],in_data[1795],in_data[1699],in_data[1603],in_data[1507],in_data[1411],in_data[1315],in_data[1219],in_data[1123],in_data[1027],in_data[931],in_data[835],in_data[739],in_data[643],in_data[547],in_data[451],in_data[355],in_data[259],in_data[163],in_data[67],in_data[12258],in_data[12162],in_data[12066],in_data[11970],in_data[11874],in_data[11778],in_data[11682],in_data[11586],in_data[11490],in_data[11394],in_data[11298],in_data[11202],in_data[11106],in_data[11010],in_data[10914],in_data[10818],in_data[10722],in_data[10626],in_data[10530],in_data[10434],in_data[10338],in_data[10242],in_data[10146],in_data[10050],in_data[9954],in_data[9858],in_data[9762],in_data[9666],in_data[9570],in_data[9474],in_data[9378],in_data[9282],in_data[9186],in_data[9090],in_data[8994],in_data[8898],in_data[8802],in_data[8706],in_data[8610],in_data[8514],in_data[8418],in_data[8322],in_data[8226],in_data[8130],in_data[8034],in_data[7938],in_data[7842],in_data[7746],in_data[7650],in_data[7554],in_data[7458],in_data[7362],in_data[7266],in_data[7170],in_data[7074],in_data[6978],in_data[6882],in_data[6786],in_data[6690],in_data[6594],in_data[6498],in_data[6402],in_data[6306],in_data[6210],in_data[6114],in_data[6018],in_data[5922],in_data[5826],in_data[5730],in_data[5634],in_data[5538],in_data[5442],in_data[5346],in_data[5250],in_data[5154],in_data[5058],in_data[4962],in_data[4866],in_data[4770],in_data[4674],in_data[4578],in_data[4482],in_data[4386],in_data[4290],in_data[4194],in_data[4098],in_data[4002],in_data[3906],in_data[3810],in_data[3714],in_data[3618],in_data[3522],in_data[3426],in_data[3330],in_data[3234],in_data[3138],in_data[3042],in_data[2946],in_data[2850],in_data[2754],in_data[2658],in_data[2562],in_data[2466],in_data[2370],in_data[2274],in_data[2178],in_data[2082],in_data[1986],in_data[1890],in_data[1794],in_data[1698],in_data[1602],in_data[1506],in_data[1410],in_data[1314],in_data[1218],in_data[1122],in_data[1026],in_data[930],in_data[834],in_data[738],in_data[642],in_data[546],in_data[450],in_data[354],in_data[258],in_data[162],in_data[66],in_data[12257],in_data[12161],in_data[12065],in_data[11969],in_data[11873],in_data[11777],in_data[11681],in_data[11585],in_data[11489],in_data[11393],in_data[11297],in_data[11201],in_data[11105],in_data[11009],in_data[10913],in_data[10817],in_data[10721],in_data[10625],in_data[10529],in_data[10433],in_data[10337],in_data[10241],in_data[10145],in_data[10049],in_data[9953],in_data[9857],in_data[9761],in_data[9665],in_data[9569],in_data[9473],in_data[9377],in_data[9281],in_data[9185],in_data[9089],in_data[8993],in_data[8897],in_data[8801],in_data[8705],in_data[8609],in_data[8513],in_data[8417],in_data[8321],in_data[8225],in_data[8129],in_data[8033],in_data[7937],in_data[7841],in_data[7745],in_data[7649],in_data[7553],in_data[7457],in_data[7361],in_data[7265],in_data[7169],in_data[7073],in_data[6977],in_data[6881],in_data[6785],in_data[6689],in_data[6593],in_data[6497],in_data[6401],in_data[6305],in_data[6209],in_data[6113],in_data[6017],in_data[5921],in_data[5825],in_data[5729],in_data[5633],in_data[5537],in_data[5441],in_data[5345],in_data[5249],in_data[5153],in_data[5057],in_data[4961],in_data[4865],in_data[4769],in_data[4673],in_data[4577],in_data[4481],in_data[4385],in_data[4289],in_data[4193],in_data[4097],in_data[4001],in_data[3905],in_data[3809],in_data[3713],in_data[3617],in_data[3521],in_data[3425],in_data[3329],in_data[3233],in_data[3137],in_data[3041],in_data[2945],in_data[2849],in_data[2753],in_data[2657],in_data[2561],in_data[2465],in_data[2369],in_data[2273],in_data[2177],in_data[2081],in_data[1985],in_data[1889],in_data[1793],in_data[1697],in_data[1601],in_data[1505],in_data[1409],in_data[1313],in_data[1217],in_data[1121],in_data[1025],in_data[929],in_data[833],in_data[737],in_data[641],in_data[545],in_data[449],in_data[353],in_data[257],in_data[161],in_data[65],in_data[12256],in_data[12160],in_data[12064],in_data[11968],in_data[11872],in_data[11776],in_data[11680],in_data[11584],in_data[11488],in_data[11392],in_data[11296],in_data[11200],in_data[11104],in_data[11008],in_data[10912],in_data[10816],in_data[10720],in_data[10624],in_data[10528],in_data[10432],in_data[10336],in_data[10240],in_data[10144],in_data[10048],in_data[9952],in_data[9856],in_data[9760],in_data[9664],in_data[9568],in_data[9472],in_data[9376],in_data[9280],in_data[9184],in_data[9088],in_data[8992],in_data[8896],in_data[8800],in_data[8704],in_data[8608],in_data[8512],in_data[8416],in_data[8320],in_data[8224],in_data[8128],in_data[8032],in_data[7936],in_data[7840],in_data[7744],in_data[7648],in_data[7552],in_data[7456],in_data[7360],in_data[7264],in_data[7168],in_data[7072],in_data[6976],in_data[6880],in_data[6784],in_data[6688],in_data[6592],in_data[6496],in_data[6400],in_data[6304],in_data[6208],in_data[6112],in_data[6016],in_data[5920],in_data[5824],in_data[5728],in_data[5632],in_data[5536],in_data[5440],in_data[5344],in_data[5248],in_data[5152],in_data[5056],in_data[4960],in_data[4864],in_data[4768],in_data[4672],in_data[4576],in_data[4480],in_data[4384],in_data[4288],in_data[4192],in_data[4096],in_data[4000],in_data[3904],in_data[3808],in_data[3712],in_data[3616],in_data[3520],in_data[3424],in_data[3328],in_data[3232],in_data[3136],in_data[3040],in_data[2944],in_data[2848],in_data[2752],in_data[2656],in_data[2560],in_data[2464],in_data[2368],in_data[2272],in_data[2176],in_data[2080],in_data[1984],in_data[1888],in_data[1792],in_data[1696],in_data[1600],in_data[1504],in_data[1408],in_data[1312],in_data[1216],in_data[1120],in_data[1024],in_data[928],in_data[832],in_data[736],in_data[640],in_data[544],in_data[448],in_data[352],in_data[256],in_data[160],in_data[64],in_data[12255],in_data[12159],in_data[12063],in_data[11967],in_data[11871],in_data[11775],in_data[11679],in_data[11583],in_data[11487],in_data[11391],in_data[11295],in_data[11199],in_data[11103],in_data[11007],in_data[10911],in_data[10815],in_data[10719],in_data[10623],in_data[10527],in_data[10431],in_data[10335],in_data[10239],in_data[10143],in_data[10047],in_data[9951],in_data[9855],in_data[9759],in_data[9663],in_data[9567],in_data[9471],in_data[9375],in_data[9279],in_data[9183],in_data[9087],in_data[8991],in_data[8895],in_data[8799],in_data[8703],in_data[8607],in_data[8511],in_data[8415],in_data[8319],in_data[8223],in_data[8127],in_data[8031],in_data[7935],in_data[7839],in_data[7743],in_data[7647],in_data[7551],in_data[7455],in_data[7359],in_data[7263],in_data[7167],in_data[7071],in_data[6975],in_data[6879],in_data[6783],in_data[6687],in_data[6591],in_data[6495],in_data[6399],in_data[6303],in_data[6207],in_data[6111],in_data[6015],in_data[5919],in_data[5823],in_data[5727],in_data[5631],in_data[5535],in_data[5439],in_data[5343],in_data[5247],in_data[5151],in_data[5055],in_data[4959],in_data[4863],in_data[4767],in_data[4671],in_data[4575],in_data[4479],in_data[4383],in_data[4287],in_data[4191],in_data[4095],in_data[3999],in_data[3903],in_data[3807],in_data[3711],in_data[3615],in_data[3519],in_data[3423],in_data[3327],in_data[3231],in_data[3135],in_data[3039],in_data[2943],in_data[2847],in_data[2751],in_data[2655],in_data[2559],in_data[2463],in_data[2367],in_data[2271],in_data[2175],in_data[2079],in_data[1983],in_data[1887],in_data[1791],in_data[1695],in_data[1599],in_data[1503],in_data[1407],in_data[1311],in_data[1215],in_data[1119],in_data[1023],in_data[927],in_data[831],in_data[735],in_data[639],in_data[543],in_data[447],in_data[351],in_data[255],in_data[159],in_data[63],in_data[12254],in_data[12158],in_data[12062],in_data[11966],in_data[11870],in_data[11774],in_data[11678],in_data[11582],in_data[11486],in_data[11390],in_data[11294],in_data[11198],in_data[11102],in_data[11006],in_data[10910],in_data[10814],in_data[10718],in_data[10622],in_data[10526],in_data[10430],in_data[10334],in_data[10238],in_data[10142],in_data[10046],in_data[9950],in_data[9854],in_data[9758],in_data[9662],in_data[9566],in_data[9470],in_data[9374],in_data[9278],in_data[9182],in_data[9086],in_data[8990],in_data[8894],in_data[8798],in_data[8702],in_data[8606],in_data[8510],in_data[8414],in_data[8318],in_data[8222],in_data[8126],in_data[8030],in_data[7934],in_data[7838],in_data[7742],in_data[7646],in_data[7550],in_data[7454],in_data[7358],in_data[7262],in_data[7166],in_data[7070],in_data[6974],in_data[6878],in_data[6782],in_data[6686],in_data[6590],in_data[6494],in_data[6398],in_data[6302],in_data[6206],in_data[6110],in_data[6014],in_data[5918],in_data[5822],in_data[5726],in_data[5630],in_data[5534],in_data[5438],in_data[5342],in_data[5246],in_data[5150],in_data[5054],in_data[4958],in_data[4862],in_data[4766],in_data[4670],in_data[4574],in_data[4478],in_data[4382],in_data[4286],in_data[4190],in_data[4094],in_data[3998],in_data[3902],in_data[3806],in_data[3710],in_data[3614],in_data[3518],in_data[3422],in_data[3326],in_data[3230],in_data[3134],in_data[3038],in_data[2942],in_data[2846],in_data[2750],in_data[2654],in_data[2558],in_data[2462],in_data[2366],in_data[2270],in_data[2174],in_data[2078],in_data[1982],in_data[1886],in_data[1790],in_data[1694],in_data[1598],in_data[1502],in_data[1406],in_data[1310],in_data[1214],in_data[1118],in_data[1022],in_data[926],in_data[830],in_data[734],in_data[638],in_data[542],in_data[446],in_data[350],in_data[254],in_data[158],in_data[62],in_data[12253],in_data[12157],in_data[12061],in_data[11965],in_data[11869],in_data[11773],in_data[11677],in_data[11581],in_data[11485],in_data[11389],in_data[11293],in_data[11197],in_data[11101],in_data[11005],in_data[10909],in_data[10813],in_data[10717],in_data[10621],in_data[10525],in_data[10429],in_data[10333],in_data[10237],in_data[10141],in_data[10045],in_data[9949],in_data[9853],in_data[9757],in_data[9661],in_data[9565],in_data[9469],in_data[9373],in_data[9277],in_data[9181],in_data[9085],in_data[8989],in_data[8893],in_data[8797],in_data[8701],in_data[8605],in_data[8509],in_data[8413],in_data[8317],in_data[8221],in_data[8125],in_data[8029],in_data[7933],in_data[7837],in_data[7741],in_data[7645],in_data[7549],in_data[7453],in_data[7357],in_data[7261],in_data[7165],in_data[7069],in_data[6973],in_data[6877],in_data[6781],in_data[6685],in_data[6589],in_data[6493],in_data[6397],in_data[6301],in_data[6205],in_data[6109],in_data[6013],in_data[5917],in_data[5821],in_data[5725],in_data[5629],in_data[5533],in_data[5437],in_data[5341],in_data[5245],in_data[5149],in_data[5053],in_data[4957],in_data[4861],in_data[4765],in_data[4669],in_data[4573],in_data[4477],in_data[4381],in_data[4285],in_data[4189],in_data[4093],in_data[3997],in_data[3901],in_data[3805],in_data[3709],in_data[3613],in_data[3517],in_data[3421],in_data[3325],in_data[3229],in_data[3133],in_data[3037],in_data[2941],in_data[2845],in_data[2749],in_data[2653],in_data[2557],in_data[2461],in_data[2365],in_data[2269],in_data[2173],in_data[2077],in_data[1981],in_data[1885],in_data[1789],in_data[1693],in_data[1597],in_data[1501],in_data[1405],in_data[1309],in_data[1213],in_data[1117],in_data[1021],in_data[925],in_data[829],in_data[733],in_data[637],in_data[541],in_data[445],in_data[349],in_data[253],in_data[157],in_data[61],in_data[12252],in_data[12156],in_data[12060],in_data[11964],in_data[11868],in_data[11772],in_data[11676],in_data[11580],in_data[11484],in_data[11388],in_data[11292],in_data[11196],in_data[11100],in_data[11004],in_data[10908],in_data[10812],in_data[10716],in_data[10620],in_data[10524],in_data[10428],in_data[10332],in_data[10236],in_data[10140],in_data[10044],in_data[9948],in_data[9852],in_data[9756],in_data[9660],in_data[9564],in_data[9468],in_data[9372],in_data[9276],in_data[9180],in_data[9084],in_data[8988],in_data[8892],in_data[8796],in_data[8700],in_data[8604],in_data[8508],in_data[8412],in_data[8316],in_data[8220],in_data[8124],in_data[8028],in_data[7932],in_data[7836],in_data[7740],in_data[7644],in_data[7548],in_data[7452],in_data[7356],in_data[7260],in_data[7164],in_data[7068],in_data[6972],in_data[6876],in_data[6780],in_data[6684],in_data[6588],in_data[6492],in_data[6396],in_data[6300],in_data[6204],in_data[6108],in_data[6012],in_data[5916],in_data[5820],in_data[5724],in_data[5628],in_data[5532],in_data[5436],in_data[5340],in_data[5244],in_data[5148],in_data[5052],in_data[4956],in_data[4860],in_data[4764],in_data[4668],in_data[4572],in_data[4476],in_data[4380],in_data[4284],in_data[4188],in_data[4092],in_data[3996],in_data[3900],in_data[3804],in_data[3708],in_data[3612],in_data[3516],in_data[3420],in_data[3324],in_data[3228],in_data[3132],in_data[3036],in_data[2940],in_data[2844],in_data[2748],in_data[2652],in_data[2556],in_data[2460],in_data[2364],in_data[2268],in_data[2172],in_data[2076],in_data[1980],in_data[1884],in_data[1788],in_data[1692],in_data[1596],in_data[1500],in_data[1404],in_data[1308],in_data[1212],in_data[1116],in_data[1020],in_data[924],in_data[828],in_data[732],in_data[636],in_data[540],in_data[444],in_data[348],in_data[252],in_data[156],in_data[60],in_data[12251],in_data[12155],in_data[12059],in_data[11963],in_data[11867],in_data[11771],in_data[11675],in_data[11579],in_data[11483],in_data[11387],in_data[11291],in_data[11195],in_data[11099],in_data[11003],in_data[10907],in_data[10811],in_data[10715],in_data[10619],in_data[10523],in_data[10427],in_data[10331],in_data[10235],in_data[10139],in_data[10043],in_data[9947],in_data[9851],in_data[9755],in_data[9659],in_data[9563],in_data[9467],in_data[9371],in_data[9275],in_data[9179],in_data[9083],in_data[8987],in_data[8891],in_data[8795],in_data[8699],in_data[8603],in_data[8507],in_data[8411],in_data[8315],in_data[8219],in_data[8123],in_data[8027],in_data[7931],in_data[7835],in_data[7739],in_data[7643],in_data[7547],in_data[7451],in_data[7355],in_data[7259],in_data[7163],in_data[7067],in_data[6971],in_data[6875],in_data[6779],in_data[6683],in_data[6587],in_data[6491],in_data[6395],in_data[6299],in_data[6203],in_data[6107],in_data[6011],in_data[5915],in_data[5819],in_data[5723],in_data[5627],in_data[5531],in_data[5435],in_data[5339],in_data[5243],in_data[5147],in_data[5051],in_data[4955],in_data[4859],in_data[4763],in_data[4667],in_data[4571],in_data[4475],in_data[4379],in_data[4283],in_data[4187],in_data[4091],in_data[3995],in_data[3899],in_data[3803],in_data[3707],in_data[3611],in_data[3515],in_data[3419],in_data[3323],in_data[3227],in_data[3131],in_data[3035],in_data[2939],in_data[2843],in_data[2747],in_data[2651],in_data[2555],in_data[2459],in_data[2363],in_data[2267],in_data[2171],in_data[2075],in_data[1979],in_data[1883],in_data[1787],in_data[1691],in_data[1595],in_data[1499],in_data[1403],in_data[1307],in_data[1211],in_data[1115],in_data[1019],in_data[923],in_data[827],in_data[731],in_data[635],in_data[539],in_data[443],in_data[347],in_data[251],in_data[155],in_data[59],in_data[12250],in_data[12154],in_data[12058],in_data[11962],in_data[11866],in_data[11770],in_data[11674],in_data[11578],in_data[11482],in_data[11386],in_data[11290],in_data[11194],in_data[11098],in_data[11002],in_data[10906],in_data[10810],in_data[10714],in_data[10618],in_data[10522],in_data[10426],in_data[10330],in_data[10234],in_data[10138],in_data[10042],in_data[9946],in_data[9850],in_data[9754],in_data[9658],in_data[9562],in_data[9466],in_data[9370],in_data[9274],in_data[9178],in_data[9082],in_data[8986],in_data[8890],in_data[8794],in_data[8698],in_data[8602],in_data[8506],in_data[8410],in_data[8314],in_data[8218],in_data[8122],in_data[8026],in_data[7930],in_data[7834],in_data[7738],in_data[7642],in_data[7546],in_data[7450],in_data[7354],in_data[7258],in_data[7162],in_data[7066],in_data[6970],in_data[6874],in_data[6778],in_data[6682],in_data[6586],in_data[6490],in_data[6394],in_data[6298],in_data[6202],in_data[6106],in_data[6010],in_data[5914],in_data[5818],in_data[5722],in_data[5626],in_data[5530],in_data[5434],in_data[5338],in_data[5242],in_data[5146],in_data[5050],in_data[4954],in_data[4858],in_data[4762],in_data[4666],in_data[4570],in_data[4474],in_data[4378],in_data[4282],in_data[4186],in_data[4090],in_data[3994],in_data[3898],in_data[3802],in_data[3706],in_data[3610],in_data[3514],in_data[3418],in_data[3322],in_data[3226],in_data[3130],in_data[3034],in_data[2938],in_data[2842],in_data[2746],in_data[2650],in_data[2554],in_data[2458],in_data[2362],in_data[2266],in_data[2170],in_data[2074],in_data[1978],in_data[1882],in_data[1786],in_data[1690],in_data[1594],in_data[1498],in_data[1402],in_data[1306],in_data[1210],in_data[1114],in_data[1018],in_data[922],in_data[826],in_data[730],in_data[634],in_data[538],in_data[442],in_data[346],in_data[250],in_data[154],in_data[58],in_data[12249],in_data[12153],in_data[12057],in_data[11961],in_data[11865],in_data[11769],in_data[11673],in_data[11577],in_data[11481],in_data[11385],in_data[11289],in_data[11193],in_data[11097],in_data[11001],in_data[10905],in_data[10809],in_data[10713],in_data[10617],in_data[10521],in_data[10425],in_data[10329],in_data[10233],in_data[10137],in_data[10041],in_data[9945],in_data[9849],in_data[9753],in_data[9657],in_data[9561],in_data[9465],in_data[9369],in_data[9273],in_data[9177],in_data[9081],in_data[8985],in_data[8889],in_data[8793],in_data[8697],in_data[8601],in_data[8505],in_data[8409],in_data[8313],in_data[8217],in_data[8121],in_data[8025],in_data[7929],in_data[7833],in_data[7737],in_data[7641],in_data[7545],in_data[7449],in_data[7353],in_data[7257],in_data[7161],in_data[7065],in_data[6969],in_data[6873],in_data[6777],in_data[6681],in_data[6585],in_data[6489],in_data[6393],in_data[6297],in_data[6201],in_data[6105],in_data[6009],in_data[5913],in_data[5817],in_data[5721],in_data[5625],in_data[5529],in_data[5433],in_data[5337],in_data[5241],in_data[5145],in_data[5049],in_data[4953],in_data[4857],in_data[4761],in_data[4665],in_data[4569],in_data[4473],in_data[4377],in_data[4281],in_data[4185],in_data[4089],in_data[3993],in_data[3897],in_data[3801],in_data[3705],in_data[3609],in_data[3513],in_data[3417],in_data[3321],in_data[3225],in_data[3129],in_data[3033],in_data[2937],in_data[2841],in_data[2745],in_data[2649],in_data[2553],in_data[2457],in_data[2361],in_data[2265],in_data[2169],in_data[2073],in_data[1977],in_data[1881],in_data[1785],in_data[1689],in_data[1593],in_data[1497],in_data[1401],in_data[1305],in_data[1209],in_data[1113],in_data[1017],in_data[921],in_data[825],in_data[729],in_data[633],in_data[537],in_data[441],in_data[345],in_data[249],in_data[153],in_data[57],in_data[12248],in_data[12152],in_data[12056],in_data[11960],in_data[11864],in_data[11768],in_data[11672],in_data[11576],in_data[11480],in_data[11384],in_data[11288],in_data[11192],in_data[11096],in_data[11000],in_data[10904],in_data[10808],in_data[10712],in_data[10616],in_data[10520],in_data[10424],in_data[10328],in_data[10232],in_data[10136],in_data[10040],in_data[9944],in_data[9848],in_data[9752],in_data[9656],in_data[9560],in_data[9464],in_data[9368],in_data[9272],in_data[9176],in_data[9080],in_data[8984],in_data[8888],in_data[8792],in_data[8696],in_data[8600],in_data[8504],in_data[8408],in_data[8312],in_data[8216],in_data[8120],in_data[8024],in_data[7928],in_data[7832],in_data[7736],in_data[7640],in_data[7544],in_data[7448],in_data[7352],in_data[7256],in_data[7160],in_data[7064],in_data[6968],in_data[6872],in_data[6776],in_data[6680],in_data[6584],in_data[6488],in_data[6392],in_data[6296],in_data[6200],in_data[6104],in_data[6008],in_data[5912],in_data[5816],in_data[5720],in_data[5624],in_data[5528],in_data[5432],in_data[5336],in_data[5240],in_data[5144],in_data[5048],in_data[4952],in_data[4856],in_data[4760],in_data[4664],in_data[4568],in_data[4472],in_data[4376],in_data[4280],in_data[4184],in_data[4088],in_data[3992],in_data[3896],in_data[3800],in_data[3704],in_data[3608],in_data[3512],in_data[3416],in_data[3320],in_data[3224],in_data[3128],in_data[3032],in_data[2936],in_data[2840],in_data[2744],in_data[2648],in_data[2552],in_data[2456],in_data[2360],in_data[2264],in_data[2168],in_data[2072],in_data[1976],in_data[1880],in_data[1784],in_data[1688],in_data[1592],in_data[1496],in_data[1400],in_data[1304],in_data[1208],in_data[1112],in_data[1016],in_data[920],in_data[824],in_data[728],in_data[632],in_data[536],in_data[440],in_data[344],in_data[248],in_data[152],in_data[56],in_data[12247],in_data[12151],in_data[12055],in_data[11959],in_data[11863],in_data[11767],in_data[11671],in_data[11575],in_data[11479],in_data[11383],in_data[11287],in_data[11191],in_data[11095],in_data[10999],in_data[10903],in_data[10807],in_data[10711],in_data[10615],in_data[10519],in_data[10423],in_data[10327],in_data[10231],in_data[10135],in_data[10039],in_data[9943],in_data[9847],in_data[9751],in_data[9655],in_data[9559],in_data[9463],in_data[9367],in_data[9271],in_data[9175],in_data[9079],in_data[8983],in_data[8887],in_data[8791],in_data[8695],in_data[8599],in_data[8503],in_data[8407],in_data[8311],in_data[8215],in_data[8119],in_data[8023],in_data[7927],in_data[7831],in_data[7735],in_data[7639],in_data[7543],in_data[7447],in_data[7351],in_data[7255],in_data[7159],in_data[7063],in_data[6967],in_data[6871],in_data[6775],in_data[6679],in_data[6583],in_data[6487],in_data[6391],in_data[6295],in_data[6199],in_data[6103],in_data[6007],in_data[5911],in_data[5815],in_data[5719],in_data[5623],in_data[5527],in_data[5431],in_data[5335],in_data[5239],in_data[5143],in_data[5047],in_data[4951],in_data[4855],in_data[4759],in_data[4663],in_data[4567],in_data[4471],in_data[4375],in_data[4279],in_data[4183],in_data[4087],in_data[3991],in_data[3895],in_data[3799],in_data[3703],in_data[3607],in_data[3511],in_data[3415],in_data[3319],in_data[3223],in_data[3127],in_data[3031],in_data[2935],in_data[2839],in_data[2743],in_data[2647],in_data[2551],in_data[2455],in_data[2359],in_data[2263],in_data[2167],in_data[2071],in_data[1975],in_data[1879],in_data[1783],in_data[1687],in_data[1591],in_data[1495],in_data[1399],in_data[1303],in_data[1207],in_data[1111],in_data[1015],in_data[919],in_data[823],in_data[727],in_data[631],in_data[535],in_data[439],in_data[343],in_data[247],in_data[151],in_data[55],in_data[12246],in_data[12150],in_data[12054],in_data[11958],in_data[11862],in_data[11766],in_data[11670],in_data[11574],in_data[11478],in_data[11382],in_data[11286],in_data[11190],in_data[11094],in_data[10998],in_data[10902],in_data[10806],in_data[10710],in_data[10614],in_data[10518],in_data[10422],in_data[10326],in_data[10230],in_data[10134],in_data[10038],in_data[9942],in_data[9846],in_data[9750],in_data[9654],in_data[9558],in_data[9462],in_data[9366],in_data[9270],in_data[9174],in_data[9078],in_data[8982],in_data[8886],in_data[8790],in_data[8694],in_data[8598],in_data[8502],in_data[8406],in_data[8310],in_data[8214],in_data[8118],in_data[8022],in_data[7926],in_data[7830],in_data[7734],in_data[7638],in_data[7542],in_data[7446],in_data[7350],in_data[7254],in_data[7158],in_data[7062],in_data[6966],in_data[6870],in_data[6774],in_data[6678],in_data[6582],in_data[6486],in_data[6390],in_data[6294],in_data[6198],in_data[6102],in_data[6006],in_data[5910],in_data[5814],in_data[5718],in_data[5622],in_data[5526],in_data[5430],in_data[5334],in_data[5238],in_data[5142],in_data[5046],in_data[4950],in_data[4854],in_data[4758],in_data[4662],in_data[4566],in_data[4470],in_data[4374],in_data[4278],in_data[4182],in_data[4086],in_data[3990],in_data[3894],in_data[3798],in_data[3702],in_data[3606],in_data[3510],in_data[3414],in_data[3318],in_data[3222],in_data[3126],in_data[3030],in_data[2934],in_data[2838],in_data[2742],in_data[2646],in_data[2550],in_data[2454],in_data[2358],in_data[2262],in_data[2166],in_data[2070],in_data[1974],in_data[1878],in_data[1782],in_data[1686],in_data[1590],in_data[1494],in_data[1398],in_data[1302],in_data[1206],in_data[1110],in_data[1014],in_data[918],in_data[822],in_data[726],in_data[630],in_data[534],in_data[438],in_data[342],in_data[246],in_data[150],in_data[54],in_data[12245],in_data[12149],in_data[12053],in_data[11957],in_data[11861],in_data[11765],in_data[11669],in_data[11573],in_data[11477],in_data[11381],in_data[11285],in_data[11189],in_data[11093],in_data[10997],in_data[10901],in_data[10805],in_data[10709],in_data[10613],in_data[10517],in_data[10421],in_data[10325],in_data[10229],in_data[10133],in_data[10037],in_data[9941],in_data[9845],in_data[9749],in_data[9653],in_data[9557],in_data[9461],in_data[9365],in_data[9269],in_data[9173],in_data[9077],in_data[8981],in_data[8885],in_data[8789],in_data[8693],in_data[8597],in_data[8501],in_data[8405],in_data[8309],in_data[8213],in_data[8117],in_data[8021],in_data[7925],in_data[7829],in_data[7733],in_data[7637],in_data[7541],in_data[7445],in_data[7349],in_data[7253],in_data[7157],in_data[7061],in_data[6965],in_data[6869],in_data[6773],in_data[6677],in_data[6581],in_data[6485],in_data[6389],in_data[6293],in_data[6197],in_data[6101],in_data[6005],in_data[5909],in_data[5813],in_data[5717],in_data[5621],in_data[5525],in_data[5429],in_data[5333],in_data[5237],in_data[5141],in_data[5045],in_data[4949],in_data[4853],in_data[4757],in_data[4661],in_data[4565],in_data[4469],in_data[4373],in_data[4277],in_data[4181],in_data[4085],in_data[3989],in_data[3893],in_data[3797],in_data[3701],in_data[3605],in_data[3509],in_data[3413],in_data[3317],in_data[3221],in_data[3125],in_data[3029],in_data[2933],in_data[2837],in_data[2741],in_data[2645],in_data[2549],in_data[2453],in_data[2357],in_data[2261],in_data[2165],in_data[2069],in_data[1973],in_data[1877],in_data[1781],in_data[1685],in_data[1589],in_data[1493],in_data[1397],in_data[1301],in_data[1205],in_data[1109],in_data[1013],in_data[917],in_data[821],in_data[725],in_data[629],in_data[533],in_data[437],in_data[341],in_data[245],in_data[149],in_data[53],in_data[12244],in_data[12148],in_data[12052],in_data[11956],in_data[11860],in_data[11764],in_data[11668],in_data[11572],in_data[11476],in_data[11380],in_data[11284],in_data[11188],in_data[11092],in_data[10996],in_data[10900],in_data[10804],in_data[10708],in_data[10612],in_data[10516],in_data[10420],in_data[10324],in_data[10228],in_data[10132],in_data[10036],in_data[9940],in_data[9844],in_data[9748],in_data[9652],in_data[9556],in_data[9460],in_data[9364],in_data[9268],in_data[9172],in_data[9076],in_data[8980],in_data[8884],in_data[8788],in_data[8692],in_data[8596],in_data[8500],in_data[8404],in_data[8308],in_data[8212],in_data[8116],in_data[8020],in_data[7924],in_data[7828],in_data[7732],in_data[7636],in_data[7540],in_data[7444],in_data[7348],in_data[7252],in_data[7156],in_data[7060],in_data[6964],in_data[6868],in_data[6772],in_data[6676],in_data[6580],in_data[6484],in_data[6388],in_data[6292],in_data[6196],in_data[6100],in_data[6004],in_data[5908],in_data[5812],in_data[5716],in_data[5620],in_data[5524],in_data[5428],in_data[5332],in_data[5236],in_data[5140],in_data[5044],in_data[4948],in_data[4852],in_data[4756],in_data[4660],in_data[4564],in_data[4468],in_data[4372],in_data[4276],in_data[4180],in_data[4084],in_data[3988],in_data[3892],in_data[3796],in_data[3700],in_data[3604],in_data[3508],in_data[3412],in_data[3316],in_data[3220],in_data[3124],in_data[3028],in_data[2932],in_data[2836],in_data[2740],in_data[2644],in_data[2548],in_data[2452],in_data[2356],in_data[2260],in_data[2164],in_data[2068],in_data[1972],in_data[1876],in_data[1780],in_data[1684],in_data[1588],in_data[1492],in_data[1396],in_data[1300],in_data[1204],in_data[1108],in_data[1012],in_data[916],in_data[820],in_data[724],in_data[628],in_data[532],in_data[436],in_data[340],in_data[244],in_data[148],in_data[52],in_data[12243],in_data[12147],in_data[12051],in_data[11955],in_data[11859],in_data[11763],in_data[11667],in_data[11571],in_data[11475],in_data[11379],in_data[11283],in_data[11187],in_data[11091],in_data[10995],in_data[10899],in_data[10803],in_data[10707],in_data[10611],in_data[10515],in_data[10419],in_data[10323],in_data[10227],in_data[10131],in_data[10035],in_data[9939],in_data[9843],in_data[9747],in_data[9651],in_data[9555],in_data[9459],in_data[9363],in_data[9267],in_data[9171],in_data[9075],in_data[8979],in_data[8883],in_data[8787],in_data[8691],in_data[8595],in_data[8499],in_data[8403],in_data[8307],in_data[8211],in_data[8115],in_data[8019],in_data[7923],in_data[7827],in_data[7731],in_data[7635],in_data[7539],in_data[7443],in_data[7347],in_data[7251],in_data[7155],in_data[7059],in_data[6963],in_data[6867],in_data[6771],in_data[6675],in_data[6579],in_data[6483],in_data[6387],in_data[6291],in_data[6195],in_data[6099],in_data[6003],in_data[5907],in_data[5811],in_data[5715],in_data[5619],in_data[5523],in_data[5427],in_data[5331],in_data[5235],in_data[5139],in_data[5043],in_data[4947],in_data[4851],in_data[4755],in_data[4659],in_data[4563],in_data[4467],in_data[4371],in_data[4275],in_data[4179],in_data[4083],in_data[3987],in_data[3891],in_data[3795],in_data[3699],in_data[3603],in_data[3507],in_data[3411],in_data[3315],in_data[3219],in_data[3123],in_data[3027],in_data[2931],in_data[2835],in_data[2739],in_data[2643],in_data[2547],in_data[2451],in_data[2355],in_data[2259],in_data[2163],in_data[2067],in_data[1971],in_data[1875],in_data[1779],in_data[1683],in_data[1587],in_data[1491],in_data[1395],in_data[1299],in_data[1203],in_data[1107],in_data[1011],in_data[915],in_data[819],in_data[723],in_data[627],in_data[531],in_data[435],in_data[339],in_data[243],in_data[147],in_data[51],in_data[12242],in_data[12146],in_data[12050],in_data[11954],in_data[11858],in_data[11762],in_data[11666],in_data[11570],in_data[11474],in_data[11378],in_data[11282],in_data[11186],in_data[11090],in_data[10994],in_data[10898],in_data[10802],in_data[10706],in_data[10610],in_data[10514],in_data[10418],in_data[10322],in_data[10226],in_data[10130],in_data[10034],in_data[9938],in_data[9842],in_data[9746],in_data[9650],in_data[9554],in_data[9458],in_data[9362],in_data[9266],in_data[9170],in_data[9074],in_data[8978],in_data[8882],in_data[8786],in_data[8690],in_data[8594],in_data[8498],in_data[8402],in_data[8306],in_data[8210],in_data[8114],in_data[8018],in_data[7922],in_data[7826],in_data[7730],in_data[7634],in_data[7538],in_data[7442],in_data[7346],in_data[7250],in_data[7154],in_data[7058],in_data[6962],in_data[6866],in_data[6770],in_data[6674],in_data[6578],in_data[6482],in_data[6386],in_data[6290],in_data[6194],in_data[6098],in_data[6002],in_data[5906],in_data[5810],in_data[5714],in_data[5618],in_data[5522],in_data[5426],in_data[5330],in_data[5234],in_data[5138],in_data[5042],in_data[4946],in_data[4850],in_data[4754],in_data[4658],in_data[4562],in_data[4466],in_data[4370],in_data[4274],in_data[4178],in_data[4082],in_data[3986],in_data[3890],in_data[3794],in_data[3698],in_data[3602],in_data[3506],in_data[3410],in_data[3314],in_data[3218],in_data[3122],in_data[3026],in_data[2930],in_data[2834],in_data[2738],in_data[2642],in_data[2546],in_data[2450],in_data[2354],in_data[2258],in_data[2162],in_data[2066],in_data[1970],in_data[1874],in_data[1778],in_data[1682],in_data[1586],in_data[1490],in_data[1394],in_data[1298],in_data[1202],in_data[1106],in_data[1010],in_data[914],in_data[818],in_data[722],in_data[626],in_data[530],in_data[434],in_data[338],in_data[242],in_data[146],in_data[50],in_data[12241],in_data[12145],in_data[12049],in_data[11953],in_data[11857],in_data[11761],in_data[11665],in_data[11569],in_data[11473],in_data[11377],in_data[11281],in_data[11185],in_data[11089],in_data[10993],in_data[10897],in_data[10801],in_data[10705],in_data[10609],in_data[10513],in_data[10417],in_data[10321],in_data[10225],in_data[10129],in_data[10033],in_data[9937],in_data[9841],in_data[9745],in_data[9649],in_data[9553],in_data[9457],in_data[9361],in_data[9265],in_data[9169],in_data[9073],in_data[8977],in_data[8881],in_data[8785],in_data[8689],in_data[8593],in_data[8497],in_data[8401],in_data[8305],in_data[8209],in_data[8113],in_data[8017],in_data[7921],in_data[7825],in_data[7729],in_data[7633],in_data[7537],in_data[7441],in_data[7345],in_data[7249],in_data[7153],in_data[7057],in_data[6961],in_data[6865],in_data[6769],in_data[6673],in_data[6577],in_data[6481],in_data[6385],in_data[6289],in_data[6193],in_data[6097],in_data[6001],in_data[5905],in_data[5809],in_data[5713],in_data[5617],in_data[5521],in_data[5425],in_data[5329],in_data[5233],in_data[5137],in_data[5041],in_data[4945],in_data[4849],in_data[4753],in_data[4657],in_data[4561],in_data[4465],in_data[4369],in_data[4273],in_data[4177],in_data[4081],in_data[3985],in_data[3889],in_data[3793],in_data[3697],in_data[3601],in_data[3505],in_data[3409],in_data[3313],in_data[3217],in_data[3121],in_data[3025],in_data[2929],in_data[2833],in_data[2737],in_data[2641],in_data[2545],in_data[2449],in_data[2353],in_data[2257],in_data[2161],in_data[2065],in_data[1969],in_data[1873],in_data[1777],in_data[1681],in_data[1585],in_data[1489],in_data[1393],in_data[1297],in_data[1201],in_data[1105],in_data[1009],in_data[913],in_data[817],in_data[721],in_data[625],in_data[529],in_data[433],in_data[337],in_data[241],in_data[145],in_data[49],in_data[12240],in_data[12144],in_data[12048],in_data[11952],in_data[11856],in_data[11760],in_data[11664],in_data[11568],in_data[11472],in_data[11376],in_data[11280],in_data[11184],in_data[11088],in_data[10992],in_data[10896],in_data[10800],in_data[10704],in_data[10608],in_data[10512],in_data[10416],in_data[10320],in_data[10224],in_data[10128],in_data[10032],in_data[9936],in_data[9840],in_data[9744],in_data[9648],in_data[9552],in_data[9456],in_data[9360],in_data[9264],in_data[9168],in_data[9072],in_data[8976],in_data[8880],in_data[8784],in_data[8688],in_data[8592],in_data[8496],in_data[8400],in_data[8304],in_data[8208],in_data[8112],in_data[8016],in_data[7920],in_data[7824],in_data[7728],in_data[7632],in_data[7536],in_data[7440],in_data[7344],in_data[7248],in_data[7152],in_data[7056],in_data[6960],in_data[6864],in_data[6768],in_data[6672],in_data[6576],in_data[6480],in_data[6384],in_data[6288],in_data[6192],in_data[6096],in_data[6000],in_data[5904],in_data[5808],in_data[5712],in_data[5616],in_data[5520],in_data[5424],in_data[5328],in_data[5232],in_data[5136],in_data[5040],in_data[4944],in_data[4848],in_data[4752],in_data[4656],in_data[4560],in_data[4464],in_data[4368],in_data[4272],in_data[4176],in_data[4080],in_data[3984],in_data[3888],in_data[3792],in_data[3696],in_data[3600],in_data[3504],in_data[3408],in_data[3312],in_data[3216],in_data[3120],in_data[3024],in_data[2928],in_data[2832],in_data[2736],in_data[2640],in_data[2544],in_data[2448],in_data[2352],in_data[2256],in_data[2160],in_data[2064],in_data[1968],in_data[1872],in_data[1776],in_data[1680],in_data[1584],in_data[1488],in_data[1392],in_data[1296],in_data[1200],in_data[1104],in_data[1008],in_data[912],in_data[816],in_data[720],in_data[624],in_data[528],in_data[432],in_data[336],in_data[240],in_data[144],in_data[48],in_data[12239],in_data[12143],in_data[12047],in_data[11951],in_data[11855],in_data[11759],in_data[11663],in_data[11567],in_data[11471],in_data[11375],in_data[11279],in_data[11183],in_data[11087],in_data[10991],in_data[10895],in_data[10799],in_data[10703],in_data[10607],in_data[10511],in_data[10415],in_data[10319],in_data[10223],in_data[10127],in_data[10031],in_data[9935],in_data[9839],in_data[9743],in_data[9647],in_data[9551],in_data[9455],in_data[9359],in_data[9263],in_data[9167],in_data[9071],in_data[8975],in_data[8879],in_data[8783],in_data[8687],in_data[8591],in_data[8495],in_data[8399],in_data[8303],in_data[8207],in_data[8111],in_data[8015],in_data[7919],in_data[7823],in_data[7727],in_data[7631],in_data[7535],in_data[7439],in_data[7343],in_data[7247],in_data[7151],in_data[7055],in_data[6959],in_data[6863],in_data[6767],in_data[6671],in_data[6575],in_data[6479],in_data[6383],in_data[6287],in_data[6191],in_data[6095],in_data[5999],in_data[5903],in_data[5807],in_data[5711],in_data[5615],in_data[5519],in_data[5423],in_data[5327],in_data[5231],in_data[5135],in_data[5039],in_data[4943],in_data[4847],in_data[4751],in_data[4655],in_data[4559],in_data[4463],in_data[4367],in_data[4271],in_data[4175],in_data[4079],in_data[3983],in_data[3887],in_data[3791],in_data[3695],in_data[3599],in_data[3503],in_data[3407],in_data[3311],in_data[3215],in_data[3119],in_data[3023],in_data[2927],in_data[2831],in_data[2735],in_data[2639],in_data[2543],in_data[2447],in_data[2351],in_data[2255],in_data[2159],in_data[2063],in_data[1967],in_data[1871],in_data[1775],in_data[1679],in_data[1583],in_data[1487],in_data[1391],in_data[1295],in_data[1199],in_data[1103],in_data[1007],in_data[911],in_data[815],in_data[719],in_data[623],in_data[527],in_data[431],in_data[335],in_data[239],in_data[143],in_data[47],in_data[12238],in_data[12142],in_data[12046],in_data[11950],in_data[11854],in_data[11758],in_data[11662],in_data[11566],in_data[11470],in_data[11374],in_data[11278],in_data[11182],in_data[11086],in_data[10990],in_data[10894],in_data[10798],in_data[10702],in_data[10606],in_data[10510],in_data[10414],in_data[10318],in_data[10222],in_data[10126],in_data[10030],in_data[9934],in_data[9838],in_data[9742],in_data[9646],in_data[9550],in_data[9454],in_data[9358],in_data[9262],in_data[9166],in_data[9070],in_data[8974],in_data[8878],in_data[8782],in_data[8686],in_data[8590],in_data[8494],in_data[8398],in_data[8302],in_data[8206],in_data[8110],in_data[8014],in_data[7918],in_data[7822],in_data[7726],in_data[7630],in_data[7534],in_data[7438],in_data[7342],in_data[7246],in_data[7150],in_data[7054],in_data[6958],in_data[6862],in_data[6766],in_data[6670],in_data[6574],in_data[6478],in_data[6382],in_data[6286],in_data[6190],in_data[6094],in_data[5998],in_data[5902],in_data[5806],in_data[5710],in_data[5614],in_data[5518],in_data[5422],in_data[5326],in_data[5230],in_data[5134],in_data[5038],in_data[4942],in_data[4846],in_data[4750],in_data[4654],in_data[4558],in_data[4462],in_data[4366],in_data[4270],in_data[4174],in_data[4078],in_data[3982],in_data[3886],in_data[3790],in_data[3694],in_data[3598],in_data[3502],in_data[3406],in_data[3310],in_data[3214],in_data[3118],in_data[3022],in_data[2926],in_data[2830],in_data[2734],in_data[2638],in_data[2542],in_data[2446],in_data[2350],in_data[2254],in_data[2158],in_data[2062],in_data[1966],in_data[1870],in_data[1774],in_data[1678],in_data[1582],in_data[1486],in_data[1390],in_data[1294],in_data[1198],in_data[1102],in_data[1006],in_data[910],in_data[814],in_data[718],in_data[622],in_data[526],in_data[430],in_data[334],in_data[238],in_data[142],in_data[46],in_data[12237],in_data[12141],in_data[12045],in_data[11949],in_data[11853],in_data[11757],in_data[11661],in_data[11565],in_data[11469],in_data[11373],in_data[11277],in_data[11181],in_data[11085],in_data[10989],in_data[10893],in_data[10797],in_data[10701],in_data[10605],in_data[10509],in_data[10413],in_data[10317],in_data[10221],in_data[10125],in_data[10029],in_data[9933],in_data[9837],in_data[9741],in_data[9645],in_data[9549],in_data[9453],in_data[9357],in_data[9261],in_data[9165],in_data[9069],in_data[8973],in_data[8877],in_data[8781],in_data[8685],in_data[8589],in_data[8493],in_data[8397],in_data[8301],in_data[8205],in_data[8109],in_data[8013],in_data[7917],in_data[7821],in_data[7725],in_data[7629],in_data[7533],in_data[7437],in_data[7341],in_data[7245],in_data[7149],in_data[7053],in_data[6957],in_data[6861],in_data[6765],in_data[6669],in_data[6573],in_data[6477],in_data[6381],in_data[6285],in_data[6189],in_data[6093],in_data[5997],in_data[5901],in_data[5805],in_data[5709],in_data[5613],in_data[5517],in_data[5421],in_data[5325],in_data[5229],in_data[5133],in_data[5037],in_data[4941],in_data[4845],in_data[4749],in_data[4653],in_data[4557],in_data[4461],in_data[4365],in_data[4269],in_data[4173],in_data[4077],in_data[3981],in_data[3885],in_data[3789],in_data[3693],in_data[3597],in_data[3501],in_data[3405],in_data[3309],in_data[3213],in_data[3117],in_data[3021],in_data[2925],in_data[2829],in_data[2733],in_data[2637],in_data[2541],in_data[2445],in_data[2349],in_data[2253],in_data[2157],in_data[2061],in_data[1965],in_data[1869],in_data[1773],in_data[1677],in_data[1581],in_data[1485],in_data[1389],in_data[1293],in_data[1197],in_data[1101],in_data[1005],in_data[909],in_data[813],in_data[717],in_data[621],in_data[525],in_data[429],in_data[333],in_data[237],in_data[141],in_data[45],in_data[12236],in_data[12140],in_data[12044],in_data[11948],in_data[11852],in_data[11756],in_data[11660],in_data[11564],in_data[11468],in_data[11372],in_data[11276],in_data[11180],in_data[11084],in_data[10988],in_data[10892],in_data[10796],in_data[10700],in_data[10604],in_data[10508],in_data[10412],in_data[10316],in_data[10220],in_data[10124],in_data[10028],in_data[9932],in_data[9836],in_data[9740],in_data[9644],in_data[9548],in_data[9452],in_data[9356],in_data[9260],in_data[9164],in_data[9068],in_data[8972],in_data[8876],in_data[8780],in_data[8684],in_data[8588],in_data[8492],in_data[8396],in_data[8300],in_data[8204],in_data[8108],in_data[8012],in_data[7916],in_data[7820],in_data[7724],in_data[7628],in_data[7532],in_data[7436],in_data[7340],in_data[7244],in_data[7148],in_data[7052],in_data[6956],in_data[6860],in_data[6764],in_data[6668],in_data[6572],in_data[6476],in_data[6380],in_data[6284],in_data[6188],in_data[6092],in_data[5996],in_data[5900],in_data[5804],in_data[5708],in_data[5612],in_data[5516],in_data[5420],in_data[5324],in_data[5228],in_data[5132],in_data[5036],in_data[4940],in_data[4844],in_data[4748],in_data[4652],in_data[4556],in_data[4460],in_data[4364],in_data[4268],in_data[4172],in_data[4076],in_data[3980],in_data[3884],in_data[3788],in_data[3692],in_data[3596],in_data[3500],in_data[3404],in_data[3308],in_data[3212],in_data[3116],in_data[3020],in_data[2924],in_data[2828],in_data[2732],in_data[2636],in_data[2540],in_data[2444],in_data[2348],in_data[2252],in_data[2156],in_data[2060],in_data[1964],in_data[1868],in_data[1772],in_data[1676],in_data[1580],in_data[1484],in_data[1388],in_data[1292],in_data[1196],in_data[1100],in_data[1004],in_data[908],in_data[812],in_data[716],in_data[620],in_data[524],in_data[428],in_data[332],in_data[236],in_data[140],in_data[44],in_data[12235],in_data[12139],in_data[12043],in_data[11947],in_data[11851],in_data[11755],in_data[11659],in_data[11563],in_data[11467],in_data[11371],in_data[11275],in_data[11179],in_data[11083],in_data[10987],in_data[10891],in_data[10795],in_data[10699],in_data[10603],in_data[10507],in_data[10411],in_data[10315],in_data[10219],in_data[10123],in_data[10027],in_data[9931],in_data[9835],in_data[9739],in_data[9643],in_data[9547],in_data[9451],in_data[9355],in_data[9259],in_data[9163],in_data[9067],in_data[8971],in_data[8875],in_data[8779],in_data[8683],in_data[8587],in_data[8491],in_data[8395],in_data[8299],in_data[8203],in_data[8107],in_data[8011],in_data[7915],in_data[7819],in_data[7723],in_data[7627],in_data[7531],in_data[7435],in_data[7339],in_data[7243],in_data[7147],in_data[7051],in_data[6955],in_data[6859],in_data[6763],in_data[6667],in_data[6571],in_data[6475],in_data[6379],in_data[6283],in_data[6187],in_data[6091],in_data[5995],in_data[5899],in_data[5803],in_data[5707],in_data[5611],in_data[5515],in_data[5419],in_data[5323],in_data[5227],in_data[5131],in_data[5035],in_data[4939],in_data[4843],in_data[4747],in_data[4651],in_data[4555],in_data[4459],in_data[4363],in_data[4267],in_data[4171],in_data[4075],in_data[3979],in_data[3883],in_data[3787],in_data[3691],in_data[3595],in_data[3499],in_data[3403],in_data[3307],in_data[3211],in_data[3115],in_data[3019],in_data[2923],in_data[2827],in_data[2731],in_data[2635],in_data[2539],in_data[2443],in_data[2347],in_data[2251],in_data[2155],in_data[2059],in_data[1963],in_data[1867],in_data[1771],in_data[1675],in_data[1579],in_data[1483],in_data[1387],in_data[1291],in_data[1195],in_data[1099],in_data[1003],in_data[907],in_data[811],in_data[715],in_data[619],in_data[523],in_data[427],in_data[331],in_data[235],in_data[139],in_data[43],in_data[12234],in_data[12138],in_data[12042],in_data[11946],in_data[11850],in_data[11754],in_data[11658],in_data[11562],in_data[11466],in_data[11370],in_data[11274],in_data[11178],in_data[11082],in_data[10986],in_data[10890],in_data[10794],in_data[10698],in_data[10602],in_data[10506],in_data[10410],in_data[10314],in_data[10218],in_data[10122],in_data[10026],in_data[9930],in_data[9834],in_data[9738],in_data[9642],in_data[9546],in_data[9450],in_data[9354],in_data[9258],in_data[9162],in_data[9066],in_data[8970],in_data[8874],in_data[8778],in_data[8682],in_data[8586],in_data[8490],in_data[8394],in_data[8298],in_data[8202],in_data[8106],in_data[8010],in_data[7914],in_data[7818],in_data[7722],in_data[7626],in_data[7530],in_data[7434],in_data[7338],in_data[7242],in_data[7146],in_data[7050],in_data[6954],in_data[6858],in_data[6762],in_data[6666],in_data[6570],in_data[6474],in_data[6378],in_data[6282],in_data[6186],in_data[6090],in_data[5994],in_data[5898],in_data[5802],in_data[5706],in_data[5610],in_data[5514],in_data[5418],in_data[5322],in_data[5226],in_data[5130],in_data[5034],in_data[4938],in_data[4842],in_data[4746],in_data[4650],in_data[4554],in_data[4458],in_data[4362],in_data[4266],in_data[4170],in_data[4074],in_data[3978],in_data[3882],in_data[3786],in_data[3690],in_data[3594],in_data[3498],in_data[3402],in_data[3306],in_data[3210],in_data[3114],in_data[3018],in_data[2922],in_data[2826],in_data[2730],in_data[2634],in_data[2538],in_data[2442],in_data[2346],in_data[2250],in_data[2154],in_data[2058],in_data[1962],in_data[1866],in_data[1770],in_data[1674],in_data[1578],in_data[1482],in_data[1386],in_data[1290],in_data[1194],in_data[1098],in_data[1002],in_data[906],in_data[810],in_data[714],in_data[618],in_data[522],in_data[426],in_data[330],in_data[234],in_data[138],in_data[42],in_data[12233],in_data[12137],in_data[12041],in_data[11945],in_data[11849],in_data[11753],in_data[11657],in_data[11561],in_data[11465],in_data[11369],in_data[11273],in_data[11177],in_data[11081],in_data[10985],in_data[10889],in_data[10793],in_data[10697],in_data[10601],in_data[10505],in_data[10409],in_data[10313],in_data[10217],in_data[10121],in_data[10025],in_data[9929],in_data[9833],in_data[9737],in_data[9641],in_data[9545],in_data[9449],in_data[9353],in_data[9257],in_data[9161],in_data[9065],in_data[8969],in_data[8873],in_data[8777],in_data[8681],in_data[8585],in_data[8489],in_data[8393],in_data[8297],in_data[8201],in_data[8105],in_data[8009],in_data[7913],in_data[7817],in_data[7721],in_data[7625],in_data[7529],in_data[7433],in_data[7337],in_data[7241],in_data[7145],in_data[7049],in_data[6953],in_data[6857],in_data[6761],in_data[6665],in_data[6569],in_data[6473],in_data[6377],in_data[6281],in_data[6185],in_data[6089],in_data[5993],in_data[5897],in_data[5801],in_data[5705],in_data[5609],in_data[5513],in_data[5417],in_data[5321],in_data[5225],in_data[5129],in_data[5033],in_data[4937],in_data[4841],in_data[4745],in_data[4649],in_data[4553],in_data[4457],in_data[4361],in_data[4265],in_data[4169],in_data[4073],in_data[3977],in_data[3881],in_data[3785],in_data[3689],in_data[3593],in_data[3497],in_data[3401],in_data[3305],in_data[3209],in_data[3113],in_data[3017],in_data[2921],in_data[2825],in_data[2729],in_data[2633],in_data[2537],in_data[2441],in_data[2345],in_data[2249],in_data[2153],in_data[2057],in_data[1961],in_data[1865],in_data[1769],in_data[1673],in_data[1577],in_data[1481],in_data[1385],in_data[1289],in_data[1193],in_data[1097],in_data[1001],in_data[905],in_data[809],in_data[713],in_data[617],in_data[521],in_data[425],in_data[329],in_data[233],in_data[137],in_data[41],in_data[12232],in_data[12136],in_data[12040],in_data[11944],in_data[11848],in_data[11752],in_data[11656],in_data[11560],in_data[11464],in_data[11368],in_data[11272],in_data[11176],in_data[11080],in_data[10984],in_data[10888],in_data[10792],in_data[10696],in_data[10600],in_data[10504],in_data[10408],in_data[10312],in_data[10216],in_data[10120],in_data[10024],in_data[9928],in_data[9832],in_data[9736],in_data[9640],in_data[9544],in_data[9448],in_data[9352],in_data[9256],in_data[9160],in_data[9064],in_data[8968],in_data[8872],in_data[8776],in_data[8680],in_data[8584],in_data[8488],in_data[8392],in_data[8296],in_data[8200],in_data[8104],in_data[8008],in_data[7912],in_data[7816],in_data[7720],in_data[7624],in_data[7528],in_data[7432],in_data[7336],in_data[7240],in_data[7144],in_data[7048],in_data[6952],in_data[6856],in_data[6760],in_data[6664],in_data[6568],in_data[6472],in_data[6376],in_data[6280],in_data[6184],in_data[6088],in_data[5992],in_data[5896],in_data[5800],in_data[5704],in_data[5608],in_data[5512],in_data[5416],in_data[5320],in_data[5224],in_data[5128],in_data[5032],in_data[4936],in_data[4840],in_data[4744],in_data[4648],in_data[4552],in_data[4456],in_data[4360],in_data[4264],in_data[4168],in_data[4072],in_data[3976],in_data[3880],in_data[3784],in_data[3688],in_data[3592],in_data[3496],in_data[3400],in_data[3304],in_data[3208],in_data[3112],in_data[3016],in_data[2920],in_data[2824],in_data[2728],in_data[2632],in_data[2536],in_data[2440],in_data[2344],in_data[2248],in_data[2152],in_data[2056],in_data[1960],in_data[1864],in_data[1768],in_data[1672],in_data[1576],in_data[1480],in_data[1384],in_data[1288],in_data[1192],in_data[1096],in_data[1000],in_data[904],in_data[808],in_data[712],in_data[616],in_data[520],in_data[424],in_data[328],in_data[232],in_data[136],in_data[40],in_data[12231],in_data[12135],in_data[12039],in_data[11943],in_data[11847],in_data[11751],in_data[11655],in_data[11559],in_data[11463],in_data[11367],in_data[11271],in_data[11175],in_data[11079],in_data[10983],in_data[10887],in_data[10791],in_data[10695],in_data[10599],in_data[10503],in_data[10407],in_data[10311],in_data[10215],in_data[10119],in_data[10023],in_data[9927],in_data[9831],in_data[9735],in_data[9639],in_data[9543],in_data[9447],in_data[9351],in_data[9255],in_data[9159],in_data[9063],in_data[8967],in_data[8871],in_data[8775],in_data[8679],in_data[8583],in_data[8487],in_data[8391],in_data[8295],in_data[8199],in_data[8103],in_data[8007],in_data[7911],in_data[7815],in_data[7719],in_data[7623],in_data[7527],in_data[7431],in_data[7335],in_data[7239],in_data[7143],in_data[7047],in_data[6951],in_data[6855],in_data[6759],in_data[6663],in_data[6567],in_data[6471],in_data[6375],in_data[6279],in_data[6183],in_data[6087],in_data[5991],in_data[5895],in_data[5799],in_data[5703],in_data[5607],in_data[5511],in_data[5415],in_data[5319],in_data[5223],in_data[5127],in_data[5031],in_data[4935],in_data[4839],in_data[4743],in_data[4647],in_data[4551],in_data[4455],in_data[4359],in_data[4263],in_data[4167],in_data[4071],in_data[3975],in_data[3879],in_data[3783],in_data[3687],in_data[3591],in_data[3495],in_data[3399],in_data[3303],in_data[3207],in_data[3111],in_data[3015],in_data[2919],in_data[2823],in_data[2727],in_data[2631],in_data[2535],in_data[2439],in_data[2343],in_data[2247],in_data[2151],in_data[2055],in_data[1959],in_data[1863],in_data[1767],in_data[1671],in_data[1575],in_data[1479],in_data[1383],in_data[1287],in_data[1191],in_data[1095],in_data[999],in_data[903],in_data[807],in_data[711],in_data[615],in_data[519],in_data[423],in_data[327],in_data[231],in_data[135],in_data[39],in_data[12230],in_data[12134],in_data[12038],in_data[11942],in_data[11846],in_data[11750],in_data[11654],in_data[11558],in_data[11462],in_data[11366],in_data[11270],in_data[11174],in_data[11078],in_data[10982],in_data[10886],in_data[10790],in_data[10694],in_data[10598],in_data[10502],in_data[10406],in_data[10310],in_data[10214],in_data[10118],in_data[10022],in_data[9926],in_data[9830],in_data[9734],in_data[9638],in_data[9542],in_data[9446],in_data[9350],in_data[9254],in_data[9158],in_data[9062],in_data[8966],in_data[8870],in_data[8774],in_data[8678],in_data[8582],in_data[8486],in_data[8390],in_data[8294],in_data[8198],in_data[8102],in_data[8006],in_data[7910],in_data[7814],in_data[7718],in_data[7622],in_data[7526],in_data[7430],in_data[7334],in_data[7238],in_data[7142],in_data[7046],in_data[6950],in_data[6854],in_data[6758],in_data[6662],in_data[6566],in_data[6470],in_data[6374],in_data[6278],in_data[6182],in_data[6086],in_data[5990],in_data[5894],in_data[5798],in_data[5702],in_data[5606],in_data[5510],in_data[5414],in_data[5318],in_data[5222],in_data[5126],in_data[5030],in_data[4934],in_data[4838],in_data[4742],in_data[4646],in_data[4550],in_data[4454],in_data[4358],in_data[4262],in_data[4166],in_data[4070],in_data[3974],in_data[3878],in_data[3782],in_data[3686],in_data[3590],in_data[3494],in_data[3398],in_data[3302],in_data[3206],in_data[3110],in_data[3014],in_data[2918],in_data[2822],in_data[2726],in_data[2630],in_data[2534],in_data[2438],in_data[2342],in_data[2246],in_data[2150],in_data[2054],in_data[1958],in_data[1862],in_data[1766],in_data[1670],in_data[1574],in_data[1478],in_data[1382],in_data[1286],in_data[1190],in_data[1094],in_data[998],in_data[902],in_data[806],in_data[710],in_data[614],in_data[518],in_data[422],in_data[326],in_data[230],in_data[134],in_data[38],in_data[12229],in_data[12133],in_data[12037],in_data[11941],in_data[11845],in_data[11749],in_data[11653],in_data[11557],in_data[11461],in_data[11365],in_data[11269],in_data[11173],in_data[11077],in_data[10981],in_data[10885],in_data[10789],in_data[10693],in_data[10597],in_data[10501],in_data[10405],in_data[10309],in_data[10213],in_data[10117],in_data[10021],in_data[9925],in_data[9829],in_data[9733],in_data[9637],in_data[9541],in_data[9445],in_data[9349],in_data[9253],in_data[9157],in_data[9061],in_data[8965],in_data[8869],in_data[8773],in_data[8677],in_data[8581],in_data[8485],in_data[8389],in_data[8293],in_data[8197],in_data[8101],in_data[8005],in_data[7909],in_data[7813],in_data[7717],in_data[7621],in_data[7525],in_data[7429],in_data[7333],in_data[7237],in_data[7141],in_data[7045],in_data[6949],in_data[6853],in_data[6757],in_data[6661],in_data[6565],in_data[6469],in_data[6373],in_data[6277],in_data[6181],in_data[6085],in_data[5989],in_data[5893],in_data[5797],in_data[5701],in_data[5605],in_data[5509],in_data[5413],in_data[5317],in_data[5221],in_data[5125],in_data[5029],in_data[4933],in_data[4837],in_data[4741],in_data[4645],in_data[4549],in_data[4453],in_data[4357],in_data[4261],in_data[4165],in_data[4069],in_data[3973],in_data[3877],in_data[3781],in_data[3685],in_data[3589],in_data[3493],in_data[3397],in_data[3301],in_data[3205],in_data[3109],in_data[3013],in_data[2917],in_data[2821],in_data[2725],in_data[2629],in_data[2533],in_data[2437],in_data[2341],in_data[2245],in_data[2149],in_data[2053],in_data[1957],in_data[1861],in_data[1765],in_data[1669],in_data[1573],in_data[1477],in_data[1381],in_data[1285],in_data[1189],in_data[1093],in_data[997],in_data[901],in_data[805],in_data[709],in_data[613],in_data[517],in_data[421],in_data[325],in_data[229],in_data[133],in_data[37],in_data[12228],in_data[12132],in_data[12036],in_data[11940],in_data[11844],in_data[11748],in_data[11652],in_data[11556],in_data[11460],in_data[11364],in_data[11268],in_data[11172],in_data[11076],in_data[10980],in_data[10884],in_data[10788],in_data[10692],in_data[10596],in_data[10500],in_data[10404],in_data[10308],in_data[10212],in_data[10116],in_data[10020],in_data[9924],in_data[9828],in_data[9732],in_data[9636],in_data[9540],in_data[9444],in_data[9348],in_data[9252],in_data[9156],in_data[9060],in_data[8964],in_data[8868],in_data[8772],in_data[8676],in_data[8580],in_data[8484],in_data[8388],in_data[8292],in_data[8196],in_data[8100],in_data[8004],in_data[7908],in_data[7812],in_data[7716],in_data[7620],in_data[7524],in_data[7428],in_data[7332],in_data[7236],in_data[7140],in_data[7044],in_data[6948],in_data[6852],in_data[6756],in_data[6660],in_data[6564],in_data[6468],in_data[6372],in_data[6276],in_data[6180],in_data[6084],in_data[5988],in_data[5892],in_data[5796],in_data[5700],in_data[5604],in_data[5508],in_data[5412],in_data[5316],in_data[5220],in_data[5124],in_data[5028],in_data[4932],in_data[4836],in_data[4740],in_data[4644],in_data[4548],in_data[4452],in_data[4356],in_data[4260],in_data[4164],in_data[4068],in_data[3972],in_data[3876],in_data[3780],in_data[3684],in_data[3588],in_data[3492],in_data[3396],in_data[3300],in_data[3204],in_data[3108],in_data[3012],in_data[2916],in_data[2820],in_data[2724],in_data[2628],in_data[2532],in_data[2436],in_data[2340],in_data[2244],in_data[2148],in_data[2052],in_data[1956],in_data[1860],in_data[1764],in_data[1668],in_data[1572],in_data[1476],in_data[1380],in_data[1284],in_data[1188],in_data[1092],in_data[996],in_data[900],in_data[804],in_data[708],in_data[612],in_data[516],in_data[420],in_data[324],in_data[228],in_data[132],in_data[36],in_data[12227],in_data[12131],in_data[12035],in_data[11939],in_data[11843],in_data[11747],in_data[11651],in_data[11555],in_data[11459],in_data[11363],in_data[11267],in_data[11171],in_data[11075],in_data[10979],in_data[10883],in_data[10787],in_data[10691],in_data[10595],in_data[10499],in_data[10403],in_data[10307],in_data[10211],in_data[10115],in_data[10019],in_data[9923],in_data[9827],in_data[9731],in_data[9635],in_data[9539],in_data[9443],in_data[9347],in_data[9251],in_data[9155],in_data[9059],in_data[8963],in_data[8867],in_data[8771],in_data[8675],in_data[8579],in_data[8483],in_data[8387],in_data[8291],in_data[8195],in_data[8099],in_data[8003],in_data[7907],in_data[7811],in_data[7715],in_data[7619],in_data[7523],in_data[7427],in_data[7331],in_data[7235],in_data[7139],in_data[7043],in_data[6947],in_data[6851],in_data[6755],in_data[6659],in_data[6563],in_data[6467],in_data[6371],in_data[6275],in_data[6179],in_data[6083],in_data[5987],in_data[5891],in_data[5795],in_data[5699],in_data[5603],in_data[5507],in_data[5411],in_data[5315],in_data[5219],in_data[5123],in_data[5027],in_data[4931],in_data[4835],in_data[4739],in_data[4643],in_data[4547],in_data[4451],in_data[4355],in_data[4259],in_data[4163],in_data[4067],in_data[3971],in_data[3875],in_data[3779],in_data[3683],in_data[3587],in_data[3491],in_data[3395],in_data[3299],in_data[3203],in_data[3107],in_data[3011],in_data[2915],in_data[2819],in_data[2723],in_data[2627],in_data[2531],in_data[2435],in_data[2339],in_data[2243],in_data[2147],in_data[2051],in_data[1955],in_data[1859],in_data[1763],in_data[1667],in_data[1571],in_data[1475],in_data[1379],in_data[1283],in_data[1187],in_data[1091],in_data[995],in_data[899],in_data[803],in_data[707],in_data[611],in_data[515],in_data[419],in_data[323],in_data[227],in_data[131],in_data[35],in_data[12226],in_data[12130],in_data[12034],in_data[11938],in_data[11842],in_data[11746],in_data[11650],in_data[11554],in_data[11458],in_data[11362],in_data[11266],in_data[11170],in_data[11074],in_data[10978],in_data[10882],in_data[10786],in_data[10690],in_data[10594],in_data[10498],in_data[10402],in_data[10306],in_data[10210],in_data[10114],in_data[10018],in_data[9922],in_data[9826],in_data[9730],in_data[9634],in_data[9538],in_data[9442],in_data[9346],in_data[9250],in_data[9154],in_data[9058],in_data[8962],in_data[8866],in_data[8770],in_data[8674],in_data[8578],in_data[8482],in_data[8386],in_data[8290],in_data[8194],in_data[8098],in_data[8002],in_data[7906],in_data[7810],in_data[7714],in_data[7618],in_data[7522],in_data[7426],in_data[7330],in_data[7234],in_data[7138],in_data[7042],in_data[6946],in_data[6850],in_data[6754],in_data[6658],in_data[6562],in_data[6466],in_data[6370],in_data[6274],in_data[6178],in_data[6082],in_data[5986],in_data[5890],in_data[5794],in_data[5698],in_data[5602],in_data[5506],in_data[5410],in_data[5314],in_data[5218],in_data[5122],in_data[5026],in_data[4930],in_data[4834],in_data[4738],in_data[4642],in_data[4546],in_data[4450],in_data[4354],in_data[4258],in_data[4162],in_data[4066],in_data[3970],in_data[3874],in_data[3778],in_data[3682],in_data[3586],in_data[3490],in_data[3394],in_data[3298],in_data[3202],in_data[3106],in_data[3010],in_data[2914],in_data[2818],in_data[2722],in_data[2626],in_data[2530],in_data[2434],in_data[2338],in_data[2242],in_data[2146],in_data[2050],in_data[1954],in_data[1858],in_data[1762],in_data[1666],in_data[1570],in_data[1474],in_data[1378],in_data[1282],in_data[1186],in_data[1090],in_data[994],in_data[898],in_data[802],in_data[706],in_data[610],in_data[514],in_data[418],in_data[322],in_data[226],in_data[130],in_data[34],in_data[12225],in_data[12129],in_data[12033],in_data[11937],in_data[11841],in_data[11745],in_data[11649],in_data[11553],in_data[11457],in_data[11361],in_data[11265],in_data[11169],in_data[11073],in_data[10977],in_data[10881],in_data[10785],in_data[10689],in_data[10593],in_data[10497],in_data[10401],in_data[10305],in_data[10209],in_data[10113],in_data[10017],in_data[9921],in_data[9825],in_data[9729],in_data[9633],in_data[9537],in_data[9441],in_data[9345],in_data[9249],in_data[9153],in_data[9057],in_data[8961],in_data[8865],in_data[8769],in_data[8673],in_data[8577],in_data[8481],in_data[8385],in_data[8289],in_data[8193],in_data[8097],in_data[8001],in_data[7905],in_data[7809],in_data[7713],in_data[7617],in_data[7521],in_data[7425],in_data[7329],in_data[7233],in_data[7137],in_data[7041],in_data[6945],in_data[6849],in_data[6753],in_data[6657],in_data[6561],in_data[6465],in_data[6369],in_data[6273],in_data[6177],in_data[6081],in_data[5985],in_data[5889],in_data[5793],in_data[5697],in_data[5601],in_data[5505],in_data[5409],in_data[5313],in_data[5217],in_data[5121],in_data[5025],in_data[4929],in_data[4833],in_data[4737],in_data[4641],in_data[4545],in_data[4449],in_data[4353],in_data[4257],in_data[4161],in_data[4065],in_data[3969],in_data[3873],in_data[3777],in_data[3681],in_data[3585],in_data[3489],in_data[3393],in_data[3297],in_data[3201],in_data[3105],in_data[3009],in_data[2913],in_data[2817],in_data[2721],in_data[2625],in_data[2529],in_data[2433],in_data[2337],in_data[2241],in_data[2145],in_data[2049],in_data[1953],in_data[1857],in_data[1761],in_data[1665],in_data[1569],in_data[1473],in_data[1377],in_data[1281],in_data[1185],in_data[1089],in_data[993],in_data[897],in_data[801],in_data[705],in_data[609],in_data[513],in_data[417],in_data[321],in_data[225],in_data[129],in_data[33],in_data[12224],in_data[12128],in_data[12032],in_data[11936],in_data[11840],in_data[11744],in_data[11648],in_data[11552],in_data[11456],in_data[11360],in_data[11264],in_data[11168],in_data[11072],in_data[10976],in_data[10880],in_data[10784],in_data[10688],in_data[10592],in_data[10496],in_data[10400],in_data[10304],in_data[10208],in_data[10112],in_data[10016],in_data[9920],in_data[9824],in_data[9728],in_data[9632],in_data[9536],in_data[9440],in_data[9344],in_data[9248],in_data[9152],in_data[9056],in_data[8960],in_data[8864],in_data[8768],in_data[8672],in_data[8576],in_data[8480],in_data[8384],in_data[8288],in_data[8192],in_data[8096],in_data[8000],in_data[7904],in_data[7808],in_data[7712],in_data[7616],in_data[7520],in_data[7424],in_data[7328],in_data[7232],in_data[7136],in_data[7040],in_data[6944],in_data[6848],in_data[6752],in_data[6656],in_data[6560],in_data[6464],in_data[6368],in_data[6272],in_data[6176],in_data[6080],in_data[5984],in_data[5888],in_data[5792],in_data[5696],in_data[5600],in_data[5504],in_data[5408],in_data[5312],in_data[5216],in_data[5120],in_data[5024],in_data[4928],in_data[4832],in_data[4736],in_data[4640],in_data[4544],in_data[4448],in_data[4352],in_data[4256],in_data[4160],in_data[4064],in_data[3968],in_data[3872],in_data[3776],in_data[3680],in_data[3584],in_data[3488],in_data[3392],in_data[3296],in_data[3200],in_data[3104],in_data[3008],in_data[2912],in_data[2816],in_data[2720],in_data[2624],in_data[2528],in_data[2432],in_data[2336],in_data[2240],in_data[2144],in_data[2048],in_data[1952],in_data[1856],in_data[1760],in_data[1664],in_data[1568],in_data[1472],in_data[1376],in_data[1280],in_data[1184],in_data[1088],in_data[992],in_data[896],in_data[800],in_data[704],in_data[608],in_data[512],in_data[416],in_data[320],in_data[224],in_data[128],in_data[32],in_data[12223],in_data[12127],in_data[12031],in_data[11935],in_data[11839],in_data[11743],in_data[11647],in_data[11551],in_data[11455],in_data[11359],in_data[11263],in_data[11167],in_data[11071],in_data[10975],in_data[10879],in_data[10783],in_data[10687],in_data[10591],in_data[10495],in_data[10399],in_data[10303],in_data[10207],in_data[10111],in_data[10015],in_data[9919],in_data[9823],in_data[9727],in_data[9631],in_data[9535],in_data[9439],in_data[9343],in_data[9247],in_data[9151],in_data[9055],in_data[8959],in_data[8863],in_data[8767],in_data[8671],in_data[8575],in_data[8479],in_data[8383],in_data[8287],in_data[8191],in_data[8095],in_data[7999],in_data[7903],in_data[7807],in_data[7711],in_data[7615],in_data[7519],in_data[7423],in_data[7327],in_data[7231],in_data[7135],in_data[7039],in_data[6943],in_data[6847],in_data[6751],in_data[6655],in_data[6559],in_data[6463],in_data[6367],in_data[6271],in_data[6175],in_data[6079],in_data[5983],in_data[5887],in_data[5791],in_data[5695],in_data[5599],in_data[5503],in_data[5407],in_data[5311],in_data[5215],in_data[5119],in_data[5023],in_data[4927],in_data[4831],in_data[4735],in_data[4639],in_data[4543],in_data[4447],in_data[4351],in_data[4255],in_data[4159],in_data[4063],in_data[3967],in_data[3871],in_data[3775],in_data[3679],in_data[3583],in_data[3487],in_data[3391],in_data[3295],in_data[3199],in_data[3103],in_data[3007],in_data[2911],in_data[2815],in_data[2719],in_data[2623],in_data[2527],in_data[2431],in_data[2335],in_data[2239],in_data[2143],in_data[2047],in_data[1951],in_data[1855],in_data[1759],in_data[1663],in_data[1567],in_data[1471],in_data[1375],in_data[1279],in_data[1183],in_data[1087],in_data[991],in_data[895],in_data[799],in_data[703],in_data[607],in_data[511],in_data[415],in_data[319],in_data[223],in_data[127],in_data[31],in_data[12222],in_data[12126],in_data[12030],in_data[11934],in_data[11838],in_data[11742],in_data[11646],in_data[11550],in_data[11454],in_data[11358],in_data[11262],in_data[11166],in_data[11070],in_data[10974],in_data[10878],in_data[10782],in_data[10686],in_data[10590],in_data[10494],in_data[10398],in_data[10302],in_data[10206],in_data[10110],in_data[10014],in_data[9918],in_data[9822],in_data[9726],in_data[9630],in_data[9534],in_data[9438],in_data[9342],in_data[9246],in_data[9150],in_data[9054],in_data[8958],in_data[8862],in_data[8766],in_data[8670],in_data[8574],in_data[8478],in_data[8382],in_data[8286],in_data[8190],in_data[8094],in_data[7998],in_data[7902],in_data[7806],in_data[7710],in_data[7614],in_data[7518],in_data[7422],in_data[7326],in_data[7230],in_data[7134],in_data[7038],in_data[6942],in_data[6846],in_data[6750],in_data[6654],in_data[6558],in_data[6462],in_data[6366],in_data[6270],in_data[6174],in_data[6078],in_data[5982],in_data[5886],in_data[5790],in_data[5694],in_data[5598],in_data[5502],in_data[5406],in_data[5310],in_data[5214],in_data[5118],in_data[5022],in_data[4926],in_data[4830],in_data[4734],in_data[4638],in_data[4542],in_data[4446],in_data[4350],in_data[4254],in_data[4158],in_data[4062],in_data[3966],in_data[3870],in_data[3774],in_data[3678],in_data[3582],in_data[3486],in_data[3390],in_data[3294],in_data[3198],in_data[3102],in_data[3006],in_data[2910],in_data[2814],in_data[2718],in_data[2622],in_data[2526],in_data[2430],in_data[2334],in_data[2238],in_data[2142],in_data[2046],in_data[1950],in_data[1854],in_data[1758],in_data[1662],in_data[1566],in_data[1470],in_data[1374],in_data[1278],in_data[1182],in_data[1086],in_data[990],in_data[894],in_data[798],in_data[702],in_data[606],in_data[510],in_data[414],in_data[318],in_data[222],in_data[126],in_data[30],in_data[12221],in_data[12125],in_data[12029],in_data[11933],in_data[11837],in_data[11741],in_data[11645],in_data[11549],in_data[11453],in_data[11357],in_data[11261],in_data[11165],in_data[11069],in_data[10973],in_data[10877],in_data[10781],in_data[10685],in_data[10589],in_data[10493],in_data[10397],in_data[10301],in_data[10205],in_data[10109],in_data[10013],in_data[9917],in_data[9821],in_data[9725],in_data[9629],in_data[9533],in_data[9437],in_data[9341],in_data[9245],in_data[9149],in_data[9053],in_data[8957],in_data[8861],in_data[8765],in_data[8669],in_data[8573],in_data[8477],in_data[8381],in_data[8285],in_data[8189],in_data[8093],in_data[7997],in_data[7901],in_data[7805],in_data[7709],in_data[7613],in_data[7517],in_data[7421],in_data[7325],in_data[7229],in_data[7133],in_data[7037],in_data[6941],in_data[6845],in_data[6749],in_data[6653],in_data[6557],in_data[6461],in_data[6365],in_data[6269],in_data[6173],in_data[6077],in_data[5981],in_data[5885],in_data[5789],in_data[5693],in_data[5597],in_data[5501],in_data[5405],in_data[5309],in_data[5213],in_data[5117],in_data[5021],in_data[4925],in_data[4829],in_data[4733],in_data[4637],in_data[4541],in_data[4445],in_data[4349],in_data[4253],in_data[4157],in_data[4061],in_data[3965],in_data[3869],in_data[3773],in_data[3677],in_data[3581],in_data[3485],in_data[3389],in_data[3293],in_data[3197],in_data[3101],in_data[3005],in_data[2909],in_data[2813],in_data[2717],in_data[2621],in_data[2525],in_data[2429],in_data[2333],in_data[2237],in_data[2141],in_data[2045],in_data[1949],in_data[1853],in_data[1757],in_data[1661],in_data[1565],in_data[1469],in_data[1373],in_data[1277],in_data[1181],in_data[1085],in_data[989],in_data[893],in_data[797],in_data[701],in_data[605],in_data[509],in_data[413],in_data[317],in_data[221],in_data[125],in_data[29],in_data[12220],in_data[12124],in_data[12028],in_data[11932],in_data[11836],in_data[11740],in_data[11644],in_data[11548],in_data[11452],in_data[11356],in_data[11260],in_data[11164],in_data[11068],in_data[10972],in_data[10876],in_data[10780],in_data[10684],in_data[10588],in_data[10492],in_data[10396],in_data[10300],in_data[10204],in_data[10108],in_data[10012],in_data[9916],in_data[9820],in_data[9724],in_data[9628],in_data[9532],in_data[9436],in_data[9340],in_data[9244],in_data[9148],in_data[9052],in_data[8956],in_data[8860],in_data[8764],in_data[8668],in_data[8572],in_data[8476],in_data[8380],in_data[8284],in_data[8188],in_data[8092],in_data[7996],in_data[7900],in_data[7804],in_data[7708],in_data[7612],in_data[7516],in_data[7420],in_data[7324],in_data[7228],in_data[7132],in_data[7036],in_data[6940],in_data[6844],in_data[6748],in_data[6652],in_data[6556],in_data[6460],in_data[6364],in_data[6268],in_data[6172],in_data[6076],in_data[5980],in_data[5884],in_data[5788],in_data[5692],in_data[5596],in_data[5500],in_data[5404],in_data[5308],in_data[5212],in_data[5116],in_data[5020],in_data[4924],in_data[4828],in_data[4732],in_data[4636],in_data[4540],in_data[4444],in_data[4348],in_data[4252],in_data[4156],in_data[4060],in_data[3964],in_data[3868],in_data[3772],in_data[3676],in_data[3580],in_data[3484],in_data[3388],in_data[3292],in_data[3196],in_data[3100],in_data[3004],in_data[2908],in_data[2812],in_data[2716],in_data[2620],in_data[2524],in_data[2428],in_data[2332],in_data[2236],in_data[2140],in_data[2044],in_data[1948],in_data[1852],in_data[1756],in_data[1660],in_data[1564],in_data[1468],in_data[1372],in_data[1276],in_data[1180],in_data[1084],in_data[988],in_data[892],in_data[796],in_data[700],in_data[604],in_data[508],in_data[412],in_data[316],in_data[220],in_data[124],in_data[28],in_data[12219],in_data[12123],in_data[12027],in_data[11931],in_data[11835],in_data[11739],in_data[11643],in_data[11547],in_data[11451],in_data[11355],in_data[11259],in_data[11163],in_data[11067],in_data[10971],in_data[10875],in_data[10779],in_data[10683],in_data[10587],in_data[10491],in_data[10395],in_data[10299],in_data[10203],in_data[10107],in_data[10011],in_data[9915],in_data[9819],in_data[9723],in_data[9627],in_data[9531],in_data[9435],in_data[9339],in_data[9243],in_data[9147],in_data[9051],in_data[8955],in_data[8859],in_data[8763],in_data[8667],in_data[8571],in_data[8475],in_data[8379],in_data[8283],in_data[8187],in_data[8091],in_data[7995],in_data[7899],in_data[7803],in_data[7707],in_data[7611],in_data[7515],in_data[7419],in_data[7323],in_data[7227],in_data[7131],in_data[7035],in_data[6939],in_data[6843],in_data[6747],in_data[6651],in_data[6555],in_data[6459],in_data[6363],in_data[6267],in_data[6171],in_data[6075],in_data[5979],in_data[5883],in_data[5787],in_data[5691],in_data[5595],in_data[5499],in_data[5403],in_data[5307],in_data[5211],in_data[5115],in_data[5019],in_data[4923],in_data[4827],in_data[4731],in_data[4635],in_data[4539],in_data[4443],in_data[4347],in_data[4251],in_data[4155],in_data[4059],in_data[3963],in_data[3867],in_data[3771],in_data[3675],in_data[3579],in_data[3483],in_data[3387],in_data[3291],in_data[3195],in_data[3099],in_data[3003],in_data[2907],in_data[2811],in_data[2715],in_data[2619],in_data[2523],in_data[2427],in_data[2331],in_data[2235],in_data[2139],in_data[2043],in_data[1947],in_data[1851],in_data[1755],in_data[1659],in_data[1563],in_data[1467],in_data[1371],in_data[1275],in_data[1179],in_data[1083],in_data[987],in_data[891],in_data[795],in_data[699],in_data[603],in_data[507],in_data[411],in_data[315],in_data[219],in_data[123],in_data[27],in_data[12218],in_data[12122],in_data[12026],in_data[11930],in_data[11834],in_data[11738],in_data[11642],in_data[11546],in_data[11450],in_data[11354],in_data[11258],in_data[11162],in_data[11066],in_data[10970],in_data[10874],in_data[10778],in_data[10682],in_data[10586],in_data[10490],in_data[10394],in_data[10298],in_data[10202],in_data[10106],in_data[10010],in_data[9914],in_data[9818],in_data[9722],in_data[9626],in_data[9530],in_data[9434],in_data[9338],in_data[9242],in_data[9146],in_data[9050],in_data[8954],in_data[8858],in_data[8762],in_data[8666],in_data[8570],in_data[8474],in_data[8378],in_data[8282],in_data[8186],in_data[8090],in_data[7994],in_data[7898],in_data[7802],in_data[7706],in_data[7610],in_data[7514],in_data[7418],in_data[7322],in_data[7226],in_data[7130],in_data[7034],in_data[6938],in_data[6842],in_data[6746],in_data[6650],in_data[6554],in_data[6458],in_data[6362],in_data[6266],in_data[6170],in_data[6074],in_data[5978],in_data[5882],in_data[5786],in_data[5690],in_data[5594],in_data[5498],in_data[5402],in_data[5306],in_data[5210],in_data[5114],in_data[5018],in_data[4922],in_data[4826],in_data[4730],in_data[4634],in_data[4538],in_data[4442],in_data[4346],in_data[4250],in_data[4154],in_data[4058],in_data[3962],in_data[3866],in_data[3770],in_data[3674],in_data[3578],in_data[3482],in_data[3386],in_data[3290],in_data[3194],in_data[3098],in_data[3002],in_data[2906],in_data[2810],in_data[2714],in_data[2618],in_data[2522],in_data[2426],in_data[2330],in_data[2234],in_data[2138],in_data[2042],in_data[1946],in_data[1850],in_data[1754],in_data[1658],in_data[1562],in_data[1466],in_data[1370],in_data[1274],in_data[1178],in_data[1082],in_data[986],in_data[890],in_data[794],in_data[698],in_data[602],in_data[506],in_data[410],in_data[314],in_data[218],in_data[122],in_data[26],in_data[12217],in_data[12121],in_data[12025],in_data[11929],in_data[11833],in_data[11737],in_data[11641],in_data[11545],in_data[11449],in_data[11353],in_data[11257],in_data[11161],in_data[11065],in_data[10969],in_data[10873],in_data[10777],in_data[10681],in_data[10585],in_data[10489],in_data[10393],in_data[10297],in_data[10201],in_data[10105],in_data[10009],in_data[9913],in_data[9817],in_data[9721],in_data[9625],in_data[9529],in_data[9433],in_data[9337],in_data[9241],in_data[9145],in_data[9049],in_data[8953],in_data[8857],in_data[8761],in_data[8665],in_data[8569],in_data[8473],in_data[8377],in_data[8281],in_data[8185],in_data[8089],in_data[7993],in_data[7897],in_data[7801],in_data[7705],in_data[7609],in_data[7513],in_data[7417],in_data[7321],in_data[7225],in_data[7129],in_data[7033],in_data[6937],in_data[6841],in_data[6745],in_data[6649],in_data[6553],in_data[6457],in_data[6361],in_data[6265],in_data[6169],in_data[6073],in_data[5977],in_data[5881],in_data[5785],in_data[5689],in_data[5593],in_data[5497],in_data[5401],in_data[5305],in_data[5209],in_data[5113],in_data[5017],in_data[4921],in_data[4825],in_data[4729],in_data[4633],in_data[4537],in_data[4441],in_data[4345],in_data[4249],in_data[4153],in_data[4057],in_data[3961],in_data[3865],in_data[3769],in_data[3673],in_data[3577],in_data[3481],in_data[3385],in_data[3289],in_data[3193],in_data[3097],in_data[3001],in_data[2905],in_data[2809],in_data[2713],in_data[2617],in_data[2521],in_data[2425],in_data[2329],in_data[2233],in_data[2137],in_data[2041],in_data[1945],in_data[1849],in_data[1753],in_data[1657],in_data[1561],in_data[1465],in_data[1369],in_data[1273],in_data[1177],in_data[1081],in_data[985],in_data[889],in_data[793],in_data[697],in_data[601],in_data[505],in_data[409],in_data[313],in_data[217],in_data[121],in_data[25],in_data[12216],in_data[12120],in_data[12024],in_data[11928],in_data[11832],in_data[11736],in_data[11640],in_data[11544],in_data[11448],in_data[11352],in_data[11256],in_data[11160],in_data[11064],in_data[10968],in_data[10872],in_data[10776],in_data[10680],in_data[10584],in_data[10488],in_data[10392],in_data[10296],in_data[10200],in_data[10104],in_data[10008],in_data[9912],in_data[9816],in_data[9720],in_data[9624],in_data[9528],in_data[9432],in_data[9336],in_data[9240],in_data[9144],in_data[9048],in_data[8952],in_data[8856],in_data[8760],in_data[8664],in_data[8568],in_data[8472],in_data[8376],in_data[8280],in_data[8184],in_data[8088],in_data[7992],in_data[7896],in_data[7800],in_data[7704],in_data[7608],in_data[7512],in_data[7416],in_data[7320],in_data[7224],in_data[7128],in_data[7032],in_data[6936],in_data[6840],in_data[6744],in_data[6648],in_data[6552],in_data[6456],in_data[6360],in_data[6264],in_data[6168],in_data[6072],in_data[5976],in_data[5880],in_data[5784],in_data[5688],in_data[5592],in_data[5496],in_data[5400],in_data[5304],in_data[5208],in_data[5112],in_data[5016],in_data[4920],in_data[4824],in_data[4728],in_data[4632],in_data[4536],in_data[4440],in_data[4344],in_data[4248],in_data[4152],in_data[4056],in_data[3960],in_data[3864],in_data[3768],in_data[3672],in_data[3576],in_data[3480],in_data[3384],in_data[3288],in_data[3192],in_data[3096],in_data[3000],in_data[2904],in_data[2808],in_data[2712],in_data[2616],in_data[2520],in_data[2424],in_data[2328],in_data[2232],in_data[2136],in_data[2040],in_data[1944],in_data[1848],in_data[1752],in_data[1656],in_data[1560],in_data[1464],in_data[1368],in_data[1272],in_data[1176],in_data[1080],in_data[984],in_data[888],in_data[792],in_data[696],in_data[600],in_data[504],in_data[408],in_data[312],in_data[216],in_data[120],in_data[24],in_data[12215],in_data[12119],in_data[12023],in_data[11927],in_data[11831],in_data[11735],in_data[11639],in_data[11543],in_data[11447],in_data[11351],in_data[11255],in_data[11159],in_data[11063],in_data[10967],in_data[10871],in_data[10775],in_data[10679],in_data[10583],in_data[10487],in_data[10391],in_data[10295],in_data[10199],in_data[10103],in_data[10007],in_data[9911],in_data[9815],in_data[9719],in_data[9623],in_data[9527],in_data[9431],in_data[9335],in_data[9239],in_data[9143],in_data[9047],in_data[8951],in_data[8855],in_data[8759],in_data[8663],in_data[8567],in_data[8471],in_data[8375],in_data[8279],in_data[8183],in_data[8087],in_data[7991],in_data[7895],in_data[7799],in_data[7703],in_data[7607],in_data[7511],in_data[7415],in_data[7319],in_data[7223],in_data[7127],in_data[7031],in_data[6935],in_data[6839],in_data[6743],in_data[6647],in_data[6551],in_data[6455],in_data[6359],in_data[6263],in_data[6167],in_data[6071],in_data[5975],in_data[5879],in_data[5783],in_data[5687],in_data[5591],in_data[5495],in_data[5399],in_data[5303],in_data[5207],in_data[5111],in_data[5015],in_data[4919],in_data[4823],in_data[4727],in_data[4631],in_data[4535],in_data[4439],in_data[4343],in_data[4247],in_data[4151],in_data[4055],in_data[3959],in_data[3863],in_data[3767],in_data[3671],in_data[3575],in_data[3479],in_data[3383],in_data[3287],in_data[3191],in_data[3095],in_data[2999],in_data[2903],in_data[2807],in_data[2711],in_data[2615],in_data[2519],in_data[2423],in_data[2327],in_data[2231],in_data[2135],in_data[2039],in_data[1943],in_data[1847],in_data[1751],in_data[1655],in_data[1559],in_data[1463],in_data[1367],in_data[1271],in_data[1175],in_data[1079],in_data[983],in_data[887],in_data[791],in_data[695],in_data[599],in_data[503],in_data[407],in_data[311],in_data[215],in_data[119],in_data[23],in_data[12214],in_data[12118],in_data[12022],in_data[11926],in_data[11830],in_data[11734],in_data[11638],in_data[11542],in_data[11446],in_data[11350],in_data[11254],in_data[11158],in_data[11062],in_data[10966],in_data[10870],in_data[10774],in_data[10678],in_data[10582],in_data[10486],in_data[10390],in_data[10294],in_data[10198],in_data[10102],in_data[10006],in_data[9910],in_data[9814],in_data[9718],in_data[9622],in_data[9526],in_data[9430],in_data[9334],in_data[9238],in_data[9142],in_data[9046],in_data[8950],in_data[8854],in_data[8758],in_data[8662],in_data[8566],in_data[8470],in_data[8374],in_data[8278],in_data[8182],in_data[8086],in_data[7990],in_data[7894],in_data[7798],in_data[7702],in_data[7606],in_data[7510],in_data[7414],in_data[7318],in_data[7222],in_data[7126],in_data[7030],in_data[6934],in_data[6838],in_data[6742],in_data[6646],in_data[6550],in_data[6454],in_data[6358],in_data[6262],in_data[6166],in_data[6070],in_data[5974],in_data[5878],in_data[5782],in_data[5686],in_data[5590],in_data[5494],in_data[5398],in_data[5302],in_data[5206],in_data[5110],in_data[5014],in_data[4918],in_data[4822],in_data[4726],in_data[4630],in_data[4534],in_data[4438],in_data[4342],in_data[4246],in_data[4150],in_data[4054],in_data[3958],in_data[3862],in_data[3766],in_data[3670],in_data[3574],in_data[3478],in_data[3382],in_data[3286],in_data[3190],in_data[3094],in_data[2998],in_data[2902],in_data[2806],in_data[2710],in_data[2614],in_data[2518],in_data[2422],in_data[2326],in_data[2230],in_data[2134],in_data[2038],in_data[1942],in_data[1846],in_data[1750],in_data[1654],in_data[1558],in_data[1462],in_data[1366],in_data[1270],in_data[1174],in_data[1078],in_data[982],in_data[886],in_data[790],in_data[694],in_data[598],in_data[502],in_data[406],in_data[310],in_data[214],in_data[118],in_data[22],in_data[12213],in_data[12117],in_data[12021],in_data[11925],in_data[11829],in_data[11733],in_data[11637],in_data[11541],in_data[11445],in_data[11349],in_data[11253],in_data[11157],in_data[11061],in_data[10965],in_data[10869],in_data[10773],in_data[10677],in_data[10581],in_data[10485],in_data[10389],in_data[10293],in_data[10197],in_data[10101],in_data[10005],in_data[9909],in_data[9813],in_data[9717],in_data[9621],in_data[9525],in_data[9429],in_data[9333],in_data[9237],in_data[9141],in_data[9045],in_data[8949],in_data[8853],in_data[8757],in_data[8661],in_data[8565],in_data[8469],in_data[8373],in_data[8277],in_data[8181],in_data[8085],in_data[7989],in_data[7893],in_data[7797],in_data[7701],in_data[7605],in_data[7509],in_data[7413],in_data[7317],in_data[7221],in_data[7125],in_data[7029],in_data[6933],in_data[6837],in_data[6741],in_data[6645],in_data[6549],in_data[6453],in_data[6357],in_data[6261],in_data[6165],in_data[6069],in_data[5973],in_data[5877],in_data[5781],in_data[5685],in_data[5589],in_data[5493],in_data[5397],in_data[5301],in_data[5205],in_data[5109],in_data[5013],in_data[4917],in_data[4821],in_data[4725],in_data[4629],in_data[4533],in_data[4437],in_data[4341],in_data[4245],in_data[4149],in_data[4053],in_data[3957],in_data[3861],in_data[3765],in_data[3669],in_data[3573],in_data[3477],in_data[3381],in_data[3285],in_data[3189],in_data[3093],in_data[2997],in_data[2901],in_data[2805],in_data[2709],in_data[2613],in_data[2517],in_data[2421],in_data[2325],in_data[2229],in_data[2133],in_data[2037],in_data[1941],in_data[1845],in_data[1749],in_data[1653],in_data[1557],in_data[1461],in_data[1365],in_data[1269],in_data[1173],in_data[1077],in_data[981],in_data[885],in_data[789],in_data[693],in_data[597],in_data[501],in_data[405],in_data[309],in_data[213],in_data[117],in_data[21],in_data[12212],in_data[12116],in_data[12020],in_data[11924],in_data[11828],in_data[11732],in_data[11636],in_data[11540],in_data[11444],in_data[11348],in_data[11252],in_data[11156],in_data[11060],in_data[10964],in_data[10868],in_data[10772],in_data[10676],in_data[10580],in_data[10484],in_data[10388],in_data[10292],in_data[10196],in_data[10100],in_data[10004],in_data[9908],in_data[9812],in_data[9716],in_data[9620],in_data[9524],in_data[9428],in_data[9332],in_data[9236],in_data[9140],in_data[9044],in_data[8948],in_data[8852],in_data[8756],in_data[8660],in_data[8564],in_data[8468],in_data[8372],in_data[8276],in_data[8180],in_data[8084],in_data[7988],in_data[7892],in_data[7796],in_data[7700],in_data[7604],in_data[7508],in_data[7412],in_data[7316],in_data[7220],in_data[7124],in_data[7028],in_data[6932],in_data[6836],in_data[6740],in_data[6644],in_data[6548],in_data[6452],in_data[6356],in_data[6260],in_data[6164],in_data[6068],in_data[5972],in_data[5876],in_data[5780],in_data[5684],in_data[5588],in_data[5492],in_data[5396],in_data[5300],in_data[5204],in_data[5108],in_data[5012],in_data[4916],in_data[4820],in_data[4724],in_data[4628],in_data[4532],in_data[4436],in_data[4340],in_data[4244],in_data[4148],in_data[4052],in_data[3956],in_data[3860],in_data[3764],in_data[3668],in_data[3572],in_data[3476],in_data[3380],in_data[3284],in_data[3188],in_data[3092],in_data[2996],in_data[2900],in_data[2804],in_data[2708],in_data[2612],in_data[2516],in_data[2420],in_data[2324],in_data[2228],in_data[2132],in_data[2036],in_data[1940],in_data[1844],in_data[1748],in_data[1652],in_data[1556],in_data[1460],in_data[1364],in_data[1268],in_data[1172],in_data[1076],in_data[980],in_data[884],in_data[788],in_data[692],in_data[596],in_data[500],in_data[404],in_data[308],in_data[212],in_data[116],in_data[20],in_data[12211],in_data[12115],in_data[12019],in_data[11923],in_data[11827],in_data[11731],in_data[11635],in_data[11539],in_data[11443],in_data[11347],in_data[11251],in_data[11155],in_data[11059],in_data[10963],in_data[10867],in_data[10771],in_data[10675],in_data[10579],in_data[10483],in_data[10387],in_data[10291],in_data[10195],in_data[10099],in_data[10003],in_data[9907],in_data[9811],in_data[9715],in_data[9619],in_data[9523],in_data[9427],in_data[9331],in_data[9235],in_data[9139],in_data[9043],in_data[8947],in_data[8851],in_data[8755],in_data[8659],in_data[8563],in_data[8467],in_data[8371],in_data[8275],in_data[8179],in_data[8083],in_data[7987],in_data[7891],in_data[7795],in_data[7699],in_data[7603],in_data[7507],in_data[7411],in_data[7315],in_data[7219],in_data[7123],in_data[7027],in_data[6931],in_data[6835],in_data[6739],in_data[6643],in_data[6547],in_data[6451],in_data[6355],in_data[6259],in_data[6163],in_data[6067],in_data[5971],in_data[5875],in_data[5779],in_data[5683],in_data[5587],in_data[5491],in_data[5395],in_data[5299],in_data[5203],in_data[5107],in_data[5011],in_data[4915],in_data[4819],in_data[4723],in_data[4627],in_data[4531],in_data[4435],in_data[4339],in_data[4243],in_data[4147],in_data[4051],in_data[3955],in_data[3859],in_data[3763],in_data[3667],in_data[3571],in_data[3475],in_data[3379],in_data[3283],in_data[3187],in_data[3091],in_data[2995],in_data[2899],in_data[2803],in_data[2707],in_data[2611],in_data[2515],in_data[2419],in_data[2323],in_data[2227],in_data[2131],in_data[2035],in_data[1939],in_data[1843],in_data[1747],in_data[1651],in_data[1555],in_data[1459],in_data[1363],in_data[1267],in_data[1171],in_data[1075],in_data[979],in_data[883],in_data[787],in_data[691],in_data[595],in_data[499],in_data[403],in_data[307],in_data[211],in_data[115],in_data[19],in_data[12210],in_data[12114],in_data[12018],in_data[11922],in_data[11826],in_data[11730],in_data[11634],in_data[11538],in_data[11442],in_data[11346],in_data[11250],in_data[11154],in_data[11058],in_data[10962],in_data[10866],in_data[10770],in_data[10674],in_data[10578],in_data[10482],in_data[10386],in_data[10290],in_data[10194],in_data[10098],in_data[10002],in_data[9906],in_data[9810],in_data[9714],in_data[9618],in_data[9522],in_data[9426],in_data[9330],in_data[9234],in_data[9138],in_data[9042],in_data[8946],in_data[8850],in_data[8754],in_data[8658],in_data[8562],in_data[8466],in_data[8370],in_data[8274],in_data[8178],in_data[8082],in_data[7986],in_data[7890],in_data[7794],in_data[7698],in_data[7602],in_data[7506],in_data[7410],in_data[7314],in_data[7218],in_data[7122],in_data[7026],in_data[6930],in_data[6834],in_data[6738],in_data[6642],in_data[6546],in_data[6450],in_data[6354],in_data[6258],in_data[6162],in_data[6066],in_data[5970],in_data[5874],in_data[5778],in_data[5682],in_data[5586],in_data[5490],in_data[5394],in_data[5298],in_data[5202],in_data[5106],in_data[5010],in_data[4914],in_data[4818],in_data[4722],in_data[4626],in_data[4530],in_data[4434],in_data[4338],in_data[4242],in_data[4146],in_data[4050],in_data[3954],in_data[3858],in_data[3762],in_data[3666],in_data[3570],in_data[3474],in_data[3378],in_data[3282],in_data[3186],in_data[3090],in_data[2994],in_data[2898],in_data[2802],in_data[2706],in_data[2610],in_data[2514],in_data[2418],in_data[2322],in_data[2226],in_data[2130],in_data[2034],in_data[1938],in_data[1842],in_data[1746],in_data[1650],in_data[1554],in_data[1458],in_data[1362],in_data[1266],in_data[1170],in_data[1074],in_data[978],in_data[882],in_data[786],in_data[690],in_data[594],in_data[498],in_data[402],in_data[306],in_data[210],in_data[114],in_data[18],in_data[12209],in_data[12113],in_data[12017],in_data[11921],in_data[11825],in_data[11729],in_data[11633],in_data[11537],in_data[11441],in_data[11345],in_data[11249],in_data[11153],in_data[11057],in_data[10961],in_data[10865],in_data[10769],in_data[10673],in_data[10577],in_data[10481],in_data[10385],in_data[10289],in_data[10193],in_data[10097],in_data[10001],in_data[9905],in_data[9809],in_data[9713],in_data[9617],in_data[9521],in_data[9425],in_data[9329],in_data[9233],in_data[9137],in_data[9041],in_data[8945],in_data[8849],in_data[8753],in_data[8657],in_data[8561],in_data[8465],in_data[8369],in_data[8273],in_data[8177],in_data[8081],in_data[7985],in_data[7889],in_data[7793],in_data[7697],in_data[7601],in_data[7505],in_data[7409],in_data[7313],in_data[7217],in_data[7121],in_data[7025],in_data[6929],in_data[6833],in_data[6737],in_data[6641],in_data[6545],in_data[6449],in_data[6353],in_data[6257],in_data[6161],in_data[6065],in_data[5969],in_data[5873],in_data[5777],in_data[5681],in_data[5585],in_data[5489],in_data[5393],in_data[5297],in_data[5201],in_data[5105],in_data[5009],in_data[4913],in_data[4817],in_data[4721],in_data[4625],in_data[4529],in_data[4433],in_data[4337],in_data[4241],in_data[4145],in_data[4049],in_data[3953],in_data[3857],in_data[3761],in_data[3665],in_data[3569],in_data[3473],in_data[3377],in_data[3281],in_data[3185],in_data[3089],in_data[2993],in_data[2897],in_data[2801],in_data[2705],in_data[2609],in_data[2513],in_data[2417],in_data[2321],in_data[2225],in_data[2129],in_data[2033],in_data[1937],in_data[1841],in_data[1745],in_data[1649],in_data[1553],in_data[1457],in_data[1361],in_data[1265],in_data[1169],in_data[1073],in_data[977],in_data[881],in_data[785],in_data[689],in_data[593],in_data[497],in_data[401],in_data[305],in_data[209],in_data[113],in_data[17],in_data[12208],in_data[12112],in_data[12016],in_data[11920],in_data[11824],in_data[11728],in_data[11632],in_data[11536],in_data[11440],in_data[11344],in_data[11248],in_data[11152],in_data[11056],in_data[10960],in_data[10864],in_data[10768],in_data[10672],in_data[10576],in_data[10480],in_data[10384],in_data[10288],in_data[10192],in_data[10096],in_data[10000],in_data[9904],in_data[9808],in_data[9712],in_data[9616],in_data[9520],in_data[9424],in_data[9328],in_data[9232],in_data[9136],in_data[9040],in_data[8944],in_data[8848],in_data[8752],in_data[8656],in_data[8560],in_data[8464],in_data[8368],in_data[8272],in_data[8176],in_data[8080],in_data[7984],in_data[7888],in_data[7792],in_data[7696],in_data[7600],in_data[7504],in_data[7408],in_data[7312],in_data[7216],in_data[7120],in_data[7024],in_data[6928],in_data[6832],in_data[6736],in_data[6640],in_data[6544],in_data[6448],in_data[6352],in_data[6256],in_data[6160],in_data[6064],in_data[5968],in_data[5872],in_data[5776],in_data[5680],in_data[5584],in_data[5488],in_data[5392],in_data[5296],in_data[5200],in_data[5104],in_data[5008],in_data[4912],in_data[4816],in_data[4720],in_data[4624],in_data[4528],in_data[4432],in_data[4336],in_data[4240],in_data[4144],in_data[4048],in_data[3952],in_data[3856],in_data[3760],in_data[3664],in_data[3568],in_data[3472],in_data[3376],in_data[3280],in_data[3184],in_data[3088],in_data[2992],in_data[2896],in_data[2800],in_data[2704],in_data[2608],in_data[2512],in_data[2416],in_data[2320],in_data[2224],in_data[2128],in_data[2032],in_data[1936],in_data[1840],in_data[1744],in_data[1648],in_data[1552],in_data[1456],in_data[1360],in_data[1264],in_data[1168],in_data[1072],in_data[976],in_data[880],in_data[784],in_data[688],in_data[592],in_data[496],in_data[400],in_data[304],in_data[208],in_data[112],in_data[16],in_data[12207],in_data[12111],in_data[12015],in_data[11919],in_data[11823],in_data[11727],in_data[11631],in_data[11535],in_data[11439],in_data[11343],in_data[11247],in_data[11151],in_data[11055],in_data[10959],in_data[10863],in_data[10767],in_data[10671],in_data[10575],in_data[10479],in_data[10383],in_data[10287],in_data[10191],in_data[10095],in_data[9999],in_data[9903],in_data[9807],in_data[9711],in_data[9615],in_data[9519],in_data[9423],in_data[9327],in_data[9231],in_data[9135],in_data[9039],in_data[8943],in_data[8847],in_data[8751],in_data[8655],in_data[8559],in_data[8463],in_data[8367],in_data[8271],in_data[8175],in_data[8079],in_data[7983],in_data[7887],in_data[7791],in_data[7695],in_data[7599],in_data[7503],in_data[7407],in_data[7311],in_data[7215],in_data[7119],in_data[7023],in_data[6927],in_data[6831],in_data[6735],in_data[6639],in_data[6543],in_data[6447],in_data[6351],in_data[6255],in_data[6159],in_data[6063],in_data[5967],in_data[5871],in_data[5775],in_data[5679],in_data[5583],in_data[5487],in_data[5391],in_data[5295],in_data[5199],in_data[5103],in_data[5007],in_data[4911],in_data[4815],in_data[4719],in_data[4623],in_data[4527],in_data[4431],in_data[4335],in_data[4239],in_data[4143],in_data[4047],in_data[3951],in_data[3855],in_data[3759],in_data[3663],in_data[3567],in_data[3471],in_data[3375],in_data[3279],in_data[3183],in_data[3087],in_data[2991],in_data[2895],in_data[2799],in_data[2703],in_data[2607],in_data[2511],in_data[2415],in_data[2319],in_data[2223],in_data[2127],in_data[2031],in_data[1935],in_data[1839],in_data[1743],in_data[1647],in_data[1551],in_data[1455],in_data[1359],in_data[1263],in_data[1167],in_data[1071],in_data[975],in_data[879],in_data[783],in_data[687],in_data[591],in_data[495],in_data[399],in_data[303],in_data[207],in_data[111],in_data[15],in_data[12206],in_data[12110],in_data[12014],in_data[11918],in_data[11822],in_data[11726],in_data[11630],in_data[11534],in_data[11438],in_data[11342],in_data[11246],in_data[11150],in_data[11054],in_data[10958],in_data[10862],in_data[10766],in_data[10670],in_data[10574],in_data[10478],in_data[10382],in_data[10286],in_data[10190],in_data[10094],in_data[9998],in_data[9902],in_data[9806],in_data[9710],in_data[9614],in_data[9518],in_data[9422],in_data[9326],in_data[9230],in_data[9134],in_data[9038],in_data[8942],in_data[8846],in_data[8750],in_data[8654],in_data[8558],in_data[8462],in_data[8366],in_data[8270],in_data[8174],in_data[8078],in_data[7982],in_data[7886],in_data[7790],in_data[7694],in_data[7598],in_data[7502],in_data[7406],in_data[7310],in_data[7214],in_data[7118],in_data[7022],in_data[6926],in_data[6830],in_data[6734],in_data[6638],in_data[6542],in_data[6446],in_data[6350],in_data[6254],in_data[6158],in_data[6062],in_data[5966],in_data[5870],in_data[5774],in_data[5678],in_data[5582],in_data[5486],in_data[5390],in_data[5294],in_data[5198],in_data[5102],in_data[5006],in_data[4910],in_data[4814],in_data[4718],in_data[4622],in_data[4526],in_data[4430],in_data[4334],in_data[4238],in_data[4142],in_data[4046],in_data[3950],in_data[3854],in_data[3758],in_data[3662],in_data[3566],in_data[3470],in_data[3374],in_data[3278],in_data[3182],in_data[3086],in_data[2990],in_data[2894],in_data[2798],in_data[2702],in_data[2606],in_data[2510],in_data[2414],in_data[2318],in_data[2222],in_data[2126],in_data[2030],in_data[1934],in_data[1838],in_data[1742],in_data[1646],in_data[1550],in_data[1454],in_data[1358],in_data[1262],in_data[1166],in_data[1070],in_data[974],in_data[878],in_data[782],in_data[686],in_data[590],in_data[494],in_data[398],in_data[302],in_data[206],in_data[110],in_data[14],in_data[12205],in_data[12109],in_data[12013],in_data[11917],in_data[11821],in_data[11725],in_data[11629],in_data[11533],in_data[11437],in_data[11341],in_data[11245],in_data[11149],in_data[11053],in_data[10957],in_data[10861],in_data[10765],in_data[10669],in_data[10573],in_data[10477],in_data[10381],in_data[10285],in_data[10189],in_data[10093],in_data[9997],in_data[9901],in_data[9805],in_data[9709],in_data[9613],in_data[9517],in_data[9421],in_data[9325],in_data[9229],in_data[9133],in_data[9037],in_data[8941],in_data[8845],in_data[8749],in_data[8653],in_data[8557],in_data[8461],in_data[8365],in_data[8269],in_data[8173],in_data[8077],in_data[7981],in_data[7885],in_data[7789],in_data[7693],in_data[7597],in_data[7501],in_data[7405],in_data[7309],in_data[7213],in_data[7117],in_data[7021],in_data[6925],in_data[6829],in_data[6733],in_data[6637],in_data[6541],in_data[6445],in_data[6349],in_data[6253],in_data[6157],in_data[6061],in_data[5965],in_data[5869],in_data[5773],in_data[5677],in_data[5581],in_data[5485],in_data[5389],in_data[5293],in_data[5197],in_data[5101],in_data[5005],in_data[4909],in_data[4813],in_data[4717],in_data[4621],in_data[4525],in_data[4429],in_data[4333],in_data[4237],in_data[4141],in_data[4045],in_data[3949],in_data[3853],in_data[3757],in_data[3661],in_data[3565],in_data[3469],in_data[3373],in_data[3277],in_data[3181],in_data[3085],in_data[2989],in_data[2893],in_data[2797],in_data[2701],in_data[2605],in_data[2509],in_data[2413],in_data[2317],in_data[2221],in_data[2125],in_data[2029],in_data[1933],in_data[1837],in_data[1741],in_data[1645],in_data[1549],in_data[1453],in_data[1357],in_data[1261],in_data[1165],in_data[1069],in_data[973],in_data[877],in_data[781],in_data[685],in_data[589],in_data[493],in_data[397],in_data[301],in_data[205],in_data[109],in_data[13],in_data[12204],in_data[12108],in_data[12012],in_data[11916],in_data[11820],in_data[11724],in_data[11628],in_data[11532],in_data[11436],in_data[11340],in_data[11244],in_data[11148],in_data[11052],in_data[10956],in_data[10860],in_data[10764],in_data[10668],in_data[10572],in_data[10476],in_data[10380],in_data[10284],in_data[10188],in_data[10092],in_data[9996],in_data[9900],in_data[9804],in_data[9708],in_data[9612],in_data[9516],in_data[9420],in_data[9324],in_data[9228],in_data[9132],in_data[9036],in_data[8940],in_data[8844],in_data[8748],in_data[8652],in_data[8556],in_data[8460],in_data[8364],in_data[8268],in_data[8172],in_data[8076],in_data[7980],in_data[7884],in_data[7788],in_data[7692],in_data[7596],in_data[7500],in_data[7404],in_data[7308],in_data[7212],in_data[7116],in_data[7020],in_data[6924],in_data[6828],in_data[6732],in_data[6636],in_data[6540],in_data[6444],in_data[6348],in_data[6252],in_data[6156],in_data[6060],in_data[5964],in_data[5868],in_data[5772],in_data[5676],in_data[5580],in_data[5484],in_data[5388],in_data[5292],in_data[5196],in_data[5100],in_data[5004],in_data[4908],in_data[4812],in_data[4716],in_data[4620],in_data[4524],in_data[4428],in_data[4332],in_data[4236],in_data[4140],in_data[4044],in_data[3948],in_data[3852],in_data[3756],in_data[3660],in_data[3564],in_data[3468],in_data[3372],in_data[3276],in_data[3180],in_data[3084],in_data[2988],in_data[2892],in_data[2796],in_data[2700],in_data[2604],in_data[2508],in_data[2412],in_data[2316],in_data[2220],in_data[2124],in_data[2028],in_data[1932],in_data[1836],in_data[1740],in_data[1644],in_data[1548],in_data[1452],in_data[1356],in_data[1260],in_data[1164],in_data[1068],in_data[972],in_data[876],in_data[780],in_data[684],in_data[588],in_data[492],in_data[396],in_data[300],in_data[204],in_data[108],in_data[12],in_data[12203],in_data[12107],in_data[12011],in_data[11915],in_data[11819],in_data[11723],in_data[11627],in_data[11531],in_data[11435],in_data[11339],in_data[11243],in_data[11147],in_data[11051],in_data[10955],in_data[10859],in_data[10763],in_data[10667],in_data[10571],in_data[10475],in_data[10379],in_data[10283],in_data[10187],in_data[10091],in_data[9995],in_data[9899],in_data[9803],in_data[9707],in_data[9611],in_data[9515],in_data[9419],in_data[9323],in_data[9227],in_data[9131],in_data[9035],in_data[8939],in_data[8843],in_data[8747],in_data[8651],in_data[8555],in_data[8459],in_data[8363],in_data[8267],in_data[8171],in_data[8075],in_data[7979],in_data[7883],in_data[7787],in_data[7691],in_data[7595],in_data[7499],in_data[7403],in_data[7307],in_data[7211],in_data[7115],in_data[7019],in_data[6923],in_data[6827],in_data[6731],in_data[6635],in_data[6539],in_data[6443],in_data[6347],in_data[6251],in_data[6155],in_data[6059],in_data[5963],in_data[5867],in_data[5771],in_data[5675],in_data[5579],in_data[5483],in_data[5387],in_data[5291],in_data[5195],in_data[5099],in_data[5003],in_data[4907],in_data[4811],in_data[4715],in_data[4619],in_data[4523],in_data[4427],in_data[4331],in_data[4235],in_data[4139],in_data[4043],in_data[3947],in_data[3851],in_data[3755],in_data[3659],in_data[3563],in_data[3467],in_data[3371],in_data[3275],in_data[3179],in_data[3083],in_data[2987],in_data[2891],in_data[2795],in_data[2699],in_data[2603],in_data[2507],in_data[2411],in_data[2315],in_data[2219],in_data[2123],in_data[2027],in_data[1931],in_data[1835],in_data[1739],in_data[1643],in_data[1547],in_data[1451],in_data[1355],in_data[1259],in_data[1163],in_data[1067],in_data[971],in_data[875],in_data[779],in_data[683],in_data[587],in_data[491],in_data[395],in_data[299],in_data[203],in_data[107],in_data[11],in_data[12202],in_data[12106],in_data[12010],in_data[11914],in_data[11818],in_data[11722],in_data[11626],in_data[11530],in_data[11434],in_data[11338],in_data[11242],in_data[11146],in_data[11050],in_data[10954],in_data[10858],in_data[10762],in_data[10666],in_data[10570],in_data[10474],in_data[10378],in_data[10282],in_data[10186],in_data[10090],in_data[9994],in_data[9898],in_data[9802],in_data[9706],in_data[9610],in_data[9514],in_data[9418],in_data[9322],in_data[9226],in_data[9130],in_data[9034],in_data[8938],in_data[8842],in_data[8746],in_data[8650],in_data[8554],in_data[8458],in_data[8362],in_data[8266],in_data[8170],in_data[8074],in_data[7978],in_data[7882],in_data[7786],in_data[7690],in_data[7594],in_data[7498],in_data[7402],in_data[7306],in_data[7210],in_data[7114],in_data[7018],in_data[6922],in_data[6826],in_data[6730],in_data[6634],in_data[6538],in_data[6442],in_data[6346],in_data[6250],in_data[6154],in_data[6058],in_data[5962],in_data[5866],in_data[5770],in_data[5674],in_data[5578],in_data[5482],in_data[5386],in_data[5290],in_data[5194],in_data[5098],in_data[5002],in_data[4906],in_data[4810],in_data[4714],in_data[4618],in_data[4522],in_data[4426],in_data[4330],in_data[4234],in_data[4138],in_data[4042],in_data[3946],in_data[3850],in_data[3754],in_data[3658],in_data[3562],in_data[3466],in_data[3370],in_data[3274],in_data[3178],in_data[3082],in_data[2986],in_data[2890],in_data[2794],in_data[2698],in_data[2602],in_data[2506],in_data[2410],in_data[2314],in_data[2218],in_data[2122],in_data[2026],in_data[1930],in_data[1834],in_data[1738],in_data[1642],in_data[1546],in_data[1450],in_data[1354],in_data[1258],in_data[1162],in_data[1066],in_data[970],in_data[874],in_data[778],in_data[682],in_data[586],in_data[490],in_data[394],in_data[298],in_data[202],in_data[106],in_data[10],in_data[12201],in_data[12105],in_data[12009],in_data[11913],in_data[11817],in_data[11721],in_data[11625],in_data[11529],in_data[11433],in_data[11337],in_data[11241],in_data[11145],in_data[11049],in_data[10953],in_data[10857],in_data[10761],in_data[10665],in_data[10569],in_data[10473],in_data[10377],in_data[10281],in_data[10185],in_data[10089],in_data[9993],in_data[9897],in_data[9801],in_data[9705],in_data[9609],in_data[9513],in_data[9417],in_data[9321],in_data[9225],in_data[9129],in_data[9033],in_data[8937],in_data[8841],in_data[8745],in_data[8649],in_data[8553],in_data[8457],in_data[8361],in_data[8265],in_data[8169],in_data[8073],in_data[7977],in_data[7881],in_data[7785],in_data[7689],in_data[7593],in_data[7497],in_data[7401],in_data[7305],in_data[7209],in_data[7113],in_data[7017],in_data[6921],in_data[6825],in_data[6729],in_data[6633],in_data[6537],in_data[6441],in_data[6345],in_data[6249],in_data[6153],in_data[6057],in_data[5961],in_data[5865],in_data[5769],in_data[5673],in_data[5577],in_data[5481],in_data[5385],in_data[5289],in_data[5193],in_data[5097],in_data[5001],in_data[4905],in_data[4809],in_data[4713],in_data[4617],in_data[4521],in_data[4425],in_data[4329],in_data[4233],in_data[4137],in_data[4041],in_data[3945],in_data[3849],in_data[3753],in_data[3657],in_data[3561],in_data[3465],in_data[3369],in_data[3273],in_data[3177],in_data[3081],in_data[2985],in_data[2889],in_data[2793],in_data[2697],in_data[2601],in_data[2505],in_data[2409],in_data[2313],in_data[2217],in_data[2121],in_data[2025],in_data[1929],in_data[1833],in_data[1737],in_data[1641],in_data[1545],in_data[1449],in_data[1353],in_data[1257],in_data[1161],in_data[1065],in_data[969],in_data[873],in_data[777],in_data[681],in_data[585],in_data[489],in_data[393],in_data[297],in_data[201],in_data[105],in_data[9],in_data[12200],in_data[12104],in_data[12008],in_data[11912],in_data[11816],in_data[11720],in_data[11624],in_data[11528],in_data[11432],in_data[11336],in_data[11240],in_data[11144],in_data[11048],in_data[10952],in_data[10856],in_data[10760],in_data[10664],in_data[10568],in_data[10472],in_data[10376],in_data[10280],in_data[10184],in_data[10088],in_data[9992],in_data[9896],in_data[9800],in_data[9704],in_data[9608],in_data[9512],in_data[9416],in_data[9320],in_data[9224],in_data[9128],in_data[9032],in_data[8936],in_data[8840],in_data[8744],in_data[8648],in_data[8552],in_data[8456],in_data[8360],in_data[8264],in_data[8168],in_data[8072],in_data[7976],in_data[7880],in_data[7784],in_data[7688],in_data[7592],in_data[7496],in_data[7400],in_data[7304],in_data[7208],in_data[7112],in_data[7016],in_data[6920],in_data[6824],in_data[6728],in_data[6632],in_data[6536],in_data[6440],in_data[6344],in_data[6248],in_data[6152],in_data[6056],in_data[5960],in_data[5864],in_data[5768],in_data[5672],in_data[5576],in_data[5480],in_data[5384],in_data[5288],in_data[5192],in_data[5096],in_data[5000],in_data[4904],in_data[4808],in_data[4712],in_data[4616],in_data[4520],in_data[4424],in_data[4328],in_data[4232],in_data[4136],in_data[4040],in_data[3944],in_data[3848],in_data[3752],in_data[3656],in_data[3560],in_data[3464],in_data[3368],in_data[3272],in_data[3176],in_data[3080],in_data[2984],in_data[2888],in_data[2792],in_data[2696],in_data[2600],in_data[2504],in_data[2408],in_data[2312],in_data[2216],in_data[2120],in_data[2024],in_data[1928],in_data[1832],in_data[1736],in_data[1640],in_data[1544],in_data[1448],in_data[1352],in_data[1256],in_data[1160],in_data[1064],in_data[968],in_data[872],in_data[776],in_data[680],in_data[584],in_data[488],in_data[392],in_data[296],in_data[200],in_data[104],in_data[8],in_data[12199],in_data[12103],in_data[12007],in_data[11911],in_data[11815],in_data[11719],in_data[11623],in_data[11527],in_data[11431],in_data[11335],in_data[11239],in_data[11143],in_data[11047],in_data[10951],in_data[10855],in_data[10759],in_data[10663],in_data[10567],in_data[10471],in_data[10375],in_data[10279],in_data[10183],in_data[10087],in_data[9991],in_data[9895],in_data[9799],in_data[9703],in_data[9607],in_data[9511],in_data[9415],in_data[9319],in_data[9223],in_data[9127],in_data[9031],in_data[8935],in_data[8839],in_data[8743],in_data[8647],in_data[8551],in_data[8455],in_data[8359],in_data[8263],in_data[8167],in_data[8071],in_data[7975],in_data[7879],in_data[7783],in_data[7687],in_data[7591],in_data[7495],in_data[7399],in_data[7303],in_data[7207],in_data[7111],in_data[7015],in_data[6919],in_data[6823],in_data[6727],in_data[6631],in_data[6535],in_data[6439],in_data[6343],in_data[6247],in_data[6151],in_data[6055],in_data[5959],in_data[5863],in_data[5767],in_data[5671],in_data[5575],in_data[5479],in_data[5383],in_data[5287],in_data[5191],in_data[5095],in_data[4999],in_data[4903],in_data[4807],in_data[4711],in_data[4615],in_data[4519],in_data[4423],in_data[4327],in_data[4231],in_data[4135],in_data[4039],in_data[3943],in_data[3847],in_data[3751],in_data[3655],in_data[3559],in_data[3463],in_data[3367],in_data[3271],in_data[3175],in_data[3079],in_data[2983],in_data[2887],in_data[2791],in_data[2695],in_data[2599],in_data[2503],in_data[2407],in_data[2311],in_data[2215],in_data[2119],in_data[2023],in_data[1927],in_data[1831],in_data[1735],in_data[1639],in_data[1543],in_data[1447],in_data[1351],in_data[1255],in_data[1159],in_data[1063],in_data[967],in_data[871],in_data[775],in_data[679],in_data[583],in_data[487],in_data[391],in_data[295],in_data[199],in_data[103],in_data[7],in_data[12198],in_data[12102],in_data[12006],in_data[11910],in_data[11814],in_data[11718],in_data[11622],in_data[11526],in_data[11430],in_data[11334],in_data[11238],in_data[11142],in_data[11046],in_data[10950],in_data[10854],in_data[10758],in_data[10662],in_data[10566],in_data[10470],in_data[10374],in_data[10278],in_data[10182],in_data[10086],in_data[9990],in_data[9894],in_data[9798],in_data[9702],in_data[9606],in_data[9510],in_data[9414],in_data[9318],in_data[9222],in_data[9126],in_data[9030],in_data[8934],in_data[8838],in_data[8742],in_data[8646],in_data[8550],in_data[8454],in_data[8358],in_data[8262],in_data[8166],in_data[8070],in_data[7974],in_data[7878],in_data[7782],in_data[7686],in_data[7590],in_data[7494],in_data[7398],in_data[7302],in_data[7206],in_data[7110],in_data[7014],in_data[6918],in_data[6822],in_data[6726],in_data[6630],in_data[6534],in_data[6438],in_data[6342],in_data[6246],in_data[6150],in_data[6054],in_data[5958],in_data[5862],in_data[5766],in_data[5670],in_data[5574],in_data[5478],in_data[5382],in_data[5286],in_data[5190],in_data[5094],in_data[4998],in_data[4902],in_data[4806],in_data[4710],in_data[4614],in_data[4518],in_data[4422],in_data[4326],in_data[4230],in_data[4134],in_data[4038],in_data[3942],in_data[3846],in_data[3750],in_data[3654],in_data[3558],in_data[3462],in_data[3366],in_data[3270],in_data[3174],in_data[3078],in_data[2982],in_data[2886],in_data[2790],in_data[2694],in_data[2598],in_data[2502],in_data[2406],in_data[2310],in_data[2214],in_data[2118],in_data[2022],in_data[1926],in_data[1830],in_data[1734],in_data[1638],in_data[1542],in_data[1446],in_data[1350],in_data[1254],in_data[1158],in_data[1062],in_data[966],in_data[870],in_data[774],in_data[678],in_data[582],in_data[486],in_data[390],in_data[294],in_data[198],in_data[102],in_data[6],in_data[12197],in_data[12101],in_data[12005],in_data[11909],in_data[11813],in_data[11717],in_data[11621],in_data[11525],in_data[11429],in_data[11333],in_data[11237],in_data[11141],in_data[11045],in_data[10949],in_data[10853],in_data[10757],in_data[10661],in_data[10565],in_data[10469],in_data[10373],in_data[10277],in_data[10181],in_data[10085],in_data[9989],in_data[9893],in_data[9797],in_data[9701],in_data[9605],in_data[9509],in_data[9413],in_data[9317],in_data[9221],in_data[9125],in_data[9029],in_data[8933],in_data[8837],in_data[8741],in_data[8645],in_data[8549],in_data[8453],in_data[8357],in_data[8261],in_data[8165],in_data[8069],in_data[7973],in_data[7877],in_data[7781],in_data[7685],in_data[7589],in_data[7493],in_data[7397],in_data[7301],in_data[7205],in_data[7109],in_data[7013],in_data[6917],in_data[6821],in_data[6725],in_data[6629],in_data[6533],in_data[6437],in_data[6341],in_data[6245],in_data[6149],in_data[6053],in_data[5957],in_data[5861],in_data[5765],in_data[5669],in_data[5573],in_data[5477],in_data[5381],in_data[5285],in_data[5189],in_data[5093],in_data[4997],in_data[4901],in_data[4805],in_data[4709],in_data[4613],in_data[4517],in_data[4421],in_data[4325],in_data[4229],in_data[4133],in_data[4037],in_data[3941],in_data[3845],in_data[3749],in_data[3653],in_data[3557],in_data[3461],in_data[3365],in_data[3269],in_data[3173],in_data[3077],in_data[2981],in_data[2885],in_data[2789],in_data[2693],in_data[2597],in_data[2501],in_data[2405],in_data[2309],in_data[2213],in_data[2117],in_data[2021],in_data[1925],in_data[1829],in_data[1733],in_data[1637],in_data[1541],in_data[1445],in_data[1349],in_data[1253],in_data[1157],in_data[1061],in_data[965],in_data[869],in_data[773],in_data[677],in_data[581],in_data[485],in_data[389],in_data[293],in_data[197],in_data[101],in_data[5],in_data[12196],in_data[12100],in_data[12004],in_data[11908],in_data[11812],in_data[11716],in_data[11620],in_data[11524],in_data[11428],in_data[11332],in_data[11236],in_data[11140],in_data[11044],in_data[10948],in_data[10852],in_data[10756],in_data[10660],in_data[10564],in_data[10468],in_data[10372],in_data[10276],in_data[10180],in_data[10084],in_data[9988],in_data[9892],in_data[9796],in_data[9700],in_data[9604],in_data[9508],in_data[9412],in_data[9316],in_data[9220],in_data[9124],in_data[9028],in_data[8932],in_data[8836],in_data[8740],in_data[8644],in_data[8548],in_data[8452],in_data[8356],in_data[8260],in_data[8164],in_data[8068],in_data[7972],in_data[7876],in_data[7780],in_data[7684],in_data[7588],in_data[7492],in_data[7396],in_data[7300],in_data[7204],in_data[7108],in_data[7012],in_data[6916],in_data[6820],in_data[6724],in_data[6628],in_data[6532],in_data[6436],in_data[6340],in_data[6244],in_data[6148],in_data[6052],in_data[5956],in_data[5860],in_data[5764],in_data[5668],in_data[5572],in_data[5476],in_data[5380],in_data[5284],in_data[5188],in_data[5092],in_data[4996],in_data[4900],in_data[4804],in_data[4708],in_data[4612],in_data[4516],in_data[4420],in_data[4324],in_data[4228],in_data[4132],in_data[4036],in_data[3940],in_data[3844],in_data[3748],in_data[3652],in_data[3556],in_data[3460],in_data[3364],in_data[3268],in_data[3172],in_data[3076],in_data[2980],in_data[2884],in_data[2788],in_data[2692],in_data[2596],in_data[2500],in_data[2404],in_data[2308],in_data[2212],in_data[2116],in_data[2020],in_data[1924],in_data[1828],in_data[1732],in_data[1636],in_data[1540],in_data[1444],in_data[1348],in_data[1252],in_data[1156],in_data[1060],in_data[964],in_data[868],in_data[772],in_data[676],in_data[580],in_data[484],in_data[388],in_data[292],in_data[196],in_data[100],in_data[4],in_data[12195],in_data[12099],in_data[12003],in_data[11907],in_data[11811],in_data[11715],in_data[11619],in_data[11523],in_data[11427],in_data[11331],in_data[11235],in_data[11139],in_data[11043],in_data[10947],in_data[10851],in_data[10755],in_data[10659],in_data[10563],in_data[10467],in_data[10371],in_data[10275],in_data[10179],in_data[10083],in_data[9987],in_data[9891],in_data[9795],in_data[9699],in_data[9603],in_data[9507],in_data[9411],in_data[9315],in_data[9219],in_data[9123],in_data[9027],in_data[8931],in_data[8835],in_data[8739],in_data[8643],in_data[8547],in_data[8451],in_data[8355],in_data[8259],in_data[8163],in_data[8067],in_data[7971],in_data[7875],in_data[7779],in_data[7683],in_data[7587],in_data[7491],in_data[7395],in_data[7299],in_data[7203],in_data[7107],in_data[7011],in_data[6915],in_data[6819],in_data[6723],in_data[6627],in_data[6531],in_data[6435],in_data[6339],in_data[6243],in_data[6147],in_data[6051],in_data[5955],in_data[5859],in_data[5763],in_data[5667],in_data[5571],in_data[5475],in_data[5379],in_data[5283],in_data[5187],in_data[5091],in_data[4995],in_data[4899],in_data[4803],in_data[4707],in_data[4611],in_data[4515],in_data[4419],in_data[4323],in_data[4227],in_data[4131],in_data[4035],in_data[3939],in_data[3843],in_data[3747],in_data[3651],in_data[3555],in_data[3459],in_data[3363],in_data[3267],in_data[3171],in_data[3075],in_data[2979],in_data[2883],in_data[2787],in_data[2691],in_data[2595],in_data[2499],in_data[2403],in_data[2307],in_data[2211],in_data[2115],in_data[2019],in_data[1923],in_data[1827],in_data[1731],in_data[1635],in_data[1539],in_data[1443],in_data[1347],in_data[1251],in_data[1155],in_data[1059],in_data[963],in_data[867],in_data[771],in_data[675],in_data[579],in_data[483],in_data[387],in_data[291],in_data[195],in_data[99],in_data[3],in_data[12194],in_data[12098],in_data[12002],in_data[11906],in_data[11810],in_data[11714],in_data[11618],in_data[11522],in_data[11426],in_data[11330],in_data[11234],in_data[11138],in_data[11042],in_data[10946],in_data[10850],in_data[10754],in_data[10658],in_data[10562],in_data[10466],in_data[10370],in_data[10274],in_data[10178],in_data[10082],in_data[9986],in_data[9890],in_data[9794],in_data[9698],in_data[9602],in_data[9506],in_data[9410],in_data[9314],in_data[9218],in_data[9122],in_data[9026],in_data[8930],in_data[8834],in_data[8738],in_data[8642],in_data[8546],in_data[8450],in_data[8354],in_data[8258],in_data[8162],in_data[8066],in_data[7970],in_data[7874],in_data[7778],in_data[7682],in_data[7586],in_data[7490],in_data[7394],in_data[7298],in_data[7202],in_data[7106],in_data[7010],in_data[6914],in_data[6818],in_data[6722],in_data[6626],in_data[6530],in_data[6434],in_data[6338],in_data[6242],in_data[6146],in_data[6050],in_data[5954],in_data[5858],in_data[5762],in_data[5666],in_data[5570],in_data[5474],in_data[5378],in_data[5282],in_data[5186],in_data[5090],in_data[4994],in_data[4898],in_data[4802],in_data[4706],in_data[4610],in_data[4514],in_data[4418],in_data[4322],in_data[4226],in_data[4130],in_data[4034],in_data[3938],in_data[3842],in_data[3746],in_data[3650],in_data[3554],in_data[3458],in_data[3362],in_data[3266],in_data[3170],in_data[3074],in_data[2978],in_data[2882],in_data[2786],in_data[2690],in_data[2594],in_data[2498],in_data[2402],in_data[2306],in_data[2210],in_data[2114],in_data[2018],in_data[1922],in_data[1826],in_data[1730],in_data[1634],in_data[1538],in_data[1442],in_data[1346],in_data[1250],in_data[1154],in_data[1058],in_data[962],in_data[866],in_data[770],in_data[674],in_data[578],in_data[482],in_data[386],in_data[290],in_data[194],in_data[98],in_data[2],in_data[12193],in_data[12097],in_data[12001],in_data[11905],in_data[11809],in_data[11713],in_data[11617],in_data[11521],in_data[11425],in_data[11329],in_data[11233],in_data[11137],in_data[11041],in_data[10945],in_data[10849],in_data[10753],in_data[10657],in_data[10561],in_data[10465],in_data[10369],in_data[10273],in_data[10177],in_data[10081],in_data[9985],in_data[9889],in_data[9793],in_data[9697],in_data[9601],in_data[9505],in_data[9409],in_data[9313],in_data[9217],in_data[9121],in_data[9025],in_data[8929],in_data[8833],in_data[8737],in_data[8641],in_data[8545],in_data[8449],in_data[8353],in_data[8257],in_data[8161],in_data[8065],in_data[7969],in_data[7873],in_data[7777],in_data[7681],in_data[7585],in_data[7489],in_data[7393],in_data[7297],in_data[7201],in_data[7105],in_data[7009],in_data[6913],in_data[6817],in_data[6721],in_data[6625],in_data[6529],in_data[6433],in_data[6337],in_data[6241],in_data[6145],in_data[6049],in_data[5953],in_data[5857],in_data[5761],in_data[5665],in_data[5569],in_data[5473],in_data[5377],in_data[5281],in_data[5185],in_data[5089],in_data[4993],in_data[4897],in_data[4801],in_data[4705],in_data[4609],in_data[4513],in_data[4417],in_data[4321],in_data[4225],in_data[4129],in_data[4033],in_data[3937],in_data[3841],in_data[3745],in_data[3649],in_data[3553],in_data[3457],in_data[3361],in_data[3265],in_data[3169],in_data[3073],in_data[2977],in_data[2881],in_data[2785],in_data[2689],in_data[2593],in_data[2497],in_data[2401],in_data[2305],in_data[2209],in_data[2113],in_data[2017],in_data[1921],in_data[1825],in_data[1729],in_data[1633],in_data[1537],in_data[1441],in_data[1345],in_data[1249],in_data[1153],in_data[1057],in_data[961],in_data[865],in_data[769],in_data[673],in_data[577],in_data[481],in_data[385],in_data[289],in_data[193],in_data[97],in_data[1],in_data[12192],in_data[12096],in_data[12000],in_data[11904],in_data[11808],in_data[11712],in_data[11616],in_data[11520],in_data[11424],in_data[11328],in_data[11232],in_data[11136],in_data[11040],in_data[10944],in_data[10848],in_data[10752],in_data[10656],in_data[10560],in_data[10464],in_data[10368],in_data[10272],in_data[10176],in_data[10080],in_data[9984],in_data[9888],in_data[9792],in_data[9696],in_data[9600],in_data[9504],in_data[9408],in_data[9312],in_data[9216],in_data[9120],in_data[9024],in_data[8928],in_data[8832],in_data[8736],in_data[8640],in_data[8544],in_data[8448],in_data[8352],in_data[8256],in_data[8160],in_data[8064],in_data[7968],in_data[7872],in_data[7776],in_data[7680],in_data[7584],in_data[7488],in_data[7392],in_data[7296],in_data[7200],in_data[7104],in_data[7008],in_data[6912],in_data[6816],in_data[6720],in_data[6624],in_data[6528],in_data[6432],in_data[6336],in_data[6240],in_data[6144],in_data[6048],in_data[5952],in_data[5856],in_data[5760],in_data[5664],in_data[5568],in_data[5472],in_data[5376],in_data[5280],in_data[5184],in_data[5088],in_data[4992],in_data[4896],in_data[4800],in_data[4704],in_data[4608],in_data[4512],in_data[4416],in_data[4320],in_data[4224],in_data[4128],in_data[4032],in_data[3936],in_data[3840],in_data[3744],in_data[3648],in_data[3552],in_data[3456],in_data[3360],in_data[3264],in_data[3168],in_data[3072],in_data[2976],in_data[2880],in_data[2784],in_data[2688],in_data[2592],in_data[2496],in_data[2400],in_data[2304],in_data[2208],in_data[2112],in_data[2016],in_data[1920],in_data[1824],in_data[1728],in_data[1632],in_data[1536],in_data[1440],in_data[1344],in_data[1248],in_data[1152],in_data[1056],in_data[960],in_data[864],in_data[768],in_data[672],in_data[576],in_data[480],in_data[384],in_data[288],in_data[192],in_data[96],in_data[0]};
    //assign in_data_reorder = {in_data[127],in_data[95],in_data[63],in_data[31],in_data[126],in_data[94],in_data[62],in_data[30],in_data[125],in_data[93],in_data[61],in_data[29],in_data[124],in_data[92],in_data[60],in_data[28],in_data[123],in_data[91],in_data[59],in_data[27],in_data[122],in_data[90],in_data[58],in_data[26],in_data[121],in_data[89],in_data[57],in_data[25],in_data[120],in_data[88],in_data[56],in_data[24],in_data[119],in_data[87],in_data[55],in_data[23],in_data[118],in_data[86],in_data[54],in_data[22],in_data[117],in_data[85],in_data[53],in_data[21],in_data[116],in_data[84],in_data[52],in_data[20],in_data[115],in_data[83],in_data[51],in_data[19],in_data[114],in_data[82],in_data[50],in_data[18],in_data[113],in_data[81],in_data[49],in_data[17],in_data[112],in_data[80],in_data[48],in_data[16],in_data[111],in_data[79],in_data[47],in_data[15],in_data[110],in_data[78],in_data[46],in_data[14],in_data[109],in_data[77],in_data[45],in_data[13],in_data[108],in_data[76],in_data[44],in_data[12],in_data[107],in_data[75],in_data[43],in_data[11],in_data[106],in_data[74],in_data[42],in_data[10],in_data[105],in_data[73],in_data[41],in_data[9],in_data[104],in_data[72],in_data[40],in_data[8],in_data[103],in_data[71],in_data[39],in_data[7],in_data[102],in_data[70],in_data[38],in_data[6],in_data[101],in_data[69],in_data[37],in_data[5],in_data[100],in_data[68],in_data[36],in_data[4],in_data[99],in_data[67],in_data[35],in_data[3],in_data[98],in_data[66],in_data[34],in_data[2],in_data[97],in_data[65],in_data[33],in_data[1],in_data[96],in_data[64],in_data[32],in_data[0]};	
	genvar i;
	generate
		for(i=0; i < DATA_WIDTH; i=i+1) begin:mux_logic
		  always@(*)
		  begin
			 in_data_shifted[(i+1)*NUM_INPUT_PORTS-1:i*NUM_INPUT_PORTS] = in_data_reorder[(i+1)*NUM_INPUT_PORTS-1:i*NUM_INPUT_PORTS] >> in_sel;
		  end
		end
	endgenerate
	
	genvar j;
    generate
        for(j=0; j < DATA_WIDTH; j=j+1) begin:mux_logic1
            always@(posedge clk)
                begin
                if(rst)
                    out_data[j] <= 0;
                else
                    out_data[j] <= in_data_shifted[j*NUM_INPUT_PORTS];
                end
        end
    endgenerate	
	
    always@(posedge clk)
    begin
    if(rst)
        out_valid <= 0;
    else
        out_valid <= in_valid >> in_sel;
    end

endmodule
