/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Module: fp_abs.v
//
//	Function:
//				Evaluate the absolute value of input floating point value
//
// Dependency:
//				N/A
//
// Latency:  0 cycle

//
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module fp_abs
#(
	parameter DATA_WIDTH = 32
)
(
	input [DATA_WIDTH-1:0] in1,
	output [DATA_WIDTH-1:0] result
);
	
	assign result = {1'b0, in1[DATA_WIDTH-2:0]};

endmodule
