module Arbitration_Unit
#(
	parameter NUM_NEIGHBOR_CELLS		= 13,
	parameter NUM_PIPELINES				= 16,
	parameter CELL_ADDR_WIDTH			= 7,
	parameter CELL_ID_WIDTH				= 3,
	parameter RDADDR_ARBITER_SIZE		= 5,
	parameter RDADDR_ARBITER_BOTTOM_SIZE = 4,
	parameter RDADDR_ARBITER_MSB		= 16,
	parameter TOTAL_CELL_NUM			= 64
)
(
	input clk,
	input rst,
	input [CELL_ID_WIDTH-1:0] cellz,
	input [NUM_PIPELINES*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:0] Local_FSM_to_Cell_read_addr,
	input [NUM_PIPELINES*(NUM_NEIGHBOR_CELLS+1)-1:0] Local_enable_reading,
	
	output [NUM_PIPELINES*(NUM_NEIGHBOR_CELLS+1)-1:0] Cell_to_FSM_read_success_bit,
	output [TOTAL_CELL_NUM*CELL_ADDR_WIDTH-1:0] FSM_to_Cell_read_addr
);

wire [(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:0] FSM_to_Cell_read_addr_1_1;
wire [(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:0] FSM_to_Cell_read_addr_1_2;
wire [(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:0] FSM_to_Cell_read_addr_1_3;
wire [(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:0] FSM_to_Cell_read_addr_1_4;
wire [(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:0] FSM_to_Cell_read_addr_2_1;
wire [(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:0] FSM_to_Cell_read_addr_2_2;
wire [(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:0] FSM_to_Cell_read_addr_2_3;
wire [(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:0] FSM_to_Cell_read_addr_2_4;
wire [(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:0] FSM_to_Cell_read_addr_3_1;
wire [(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:0] FSM_to_Cell_read_addr_3_2;
wire [(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:0] FSM_to_Cell_read_addr_3_3;
wire [(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:0] FSM_to_Cell_read_addr_3_4;
wire [(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:0] FSM_to_Cell_read_addr_4_1;
wire [(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:0] FSM_to_Cell_read_addr_4_2;
wire [(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:0] FSM_to_Cell_read_addr_4_3;
wire [(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:0] FSM_to_Cell_read_addr_4_4;
assign FSM_to_Cell_read_addr_1_1 = Local_FSM_to_Cell_read_addr[1*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:0*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH];
assign FSM_to_Cell_read_addr_1_2 = Local_FSM_to_Cell_read_addr[2*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:1*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH];
assign FSM_to_Cell_read_addr_1_3 = Local_FSM_to_Cell_read_addr[3*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:2*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH];
assign FSM_to_Cell_read_addr_1_4 = Local_FSM_to_Cell_read_addr[4*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:3*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH];
assign FSM_to_Cell_read_addr_2_1 = Local_FSM_to_Cell_read_addr[5*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:4*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH];
assign FSM_to_Cell_read_addr_2_2 = Local_FSM_to_Cell_read_addr[6*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:5*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH];
assign FSM_to_Cell_read_addr_2_3 = Local_FSM_to_Cell_read_addr[7*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:6*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH];
assign FSM_to_Cell_read_addr_2_4 = Local_FSM_to_Cell_read_addr[8*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:7*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH];
assign FSM_to_Cell_read_addr_3_1 = Local_FSM_to_Cell_read_addr[9*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:8*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH];
assign FSM_to_Cell_read_addr_3_2 = Local_FSM_to_Cell_read_addr[10*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:9*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH];
assign FSM_to_Cell_read_addr_3_3 = Local_FSM_to_Cell_read_addr[11*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:10*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH];
assign FSM_to_Cell_read_addr_3_4 = Local_FSM_to_Cell_read_addr[12*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:11*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH];
assign FSM_to_Cell_read_addr_4_1 = Local_FSM_to_Cell_read_addr[13*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:12*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH];
assign FSM_to_Cell_read_addr_4_2 = Local_FSM_to_Cell_read_addr[14*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:13*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH];
assign FSM_to_Cell_read_addr_4_3 = Local_FSM_to_Cell_read_addr[15*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:14*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH];
assign FSM_to_Cell_read_addr_4_4 = Local_FSM_to_Cell_read_addr[16*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:15*(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH];

wire [NUM_NEIGHBOR_CELLS:0] enable_reading_1_1;
wire [NUM_NEIGHBOR_CELLS:0] enable_reading_1_2;
wire [NUM_NEIGHBOR_CELLS:0] enable_reading_1_3;
wire [NUM_NEIGHBOR_CELLS:0] enable_reading_1_4;
wire [NUM_NEIGHBOR_CELLS:0] enable_reading_2_1;
wire [NUM_NEIGHBOR_CELLS:0] enable_reading_2_2;
wire [NUM_NEIGHBOR_CELLS:0] enable_reading_2_3;
wire [NUM_NEIGHBOR_CELLS:0] enable_reading_2_4;
wire [NUM_NEIGHBOR_CELLS:0] enable_reading_3_1;
wire [NUM_NEIGHBOR_CELLS:0] enable_reading_3_2;
wire [NUM_NEIGHBOR_CELLS:0] enable_reading_3_3;
wire [NUM_NEIGHBOR_CELLS:0] enable_reading_3_4;
wire [NUM_NEIGHBOR_CELLS:0] enable_reading_4_1;
wire [NUM_NEIGHBOR_CELLS:0] enable_reading_4_2;
wire [NUM_NEIGHBOR_CELLS:0] enable_reading_4_3;
wire [NUM_NEIGHBOR_CELLS:0] enable_reading_4_4;
assign enable_reading_1_1 = Local_enable_reading[1*(NUM_NEIGHBOR_CELLS+1)-1:0*(NUM_NEIGHBOR_CELLS+1)];
assign enable_reading_1_2 = Local_enable_reading[2*(NUM_NEIGHBOR_CELLS+1)-1:1*(NUM_NEIGHBOR_CELLS+1)];
assign enable_reading_1_3 = Local_enable_reading[3*(NUM_NEIGHBOR_CELLS+1)-1:2*(NUM_NEIGHBOR_CELLS+1)];
assign enable_reading_1_4 = Local_enable_reading[4*(NUM_NEIGHBOR_CELLS+1)-1:3*(NUM_NEIGHBOR_CELLS+1)];
assign enable_reading_2_1 = Local_enable_reading[5*(NUM_NEIGHBOR_CELLS+1)-1:4*(NUM_NEIGHBOR_CELLS+1)];
assign enable_reading_2_2 = Local_enable_reading[6*(NUM_NEIGHBOR_CELLS+1)-1:5*(NUM_NEIGHBOR_CELLS+1)];
assign enable_reading_2_3 = Local_enable_reading[7*(NUM_NEIGHBOR_CELLS+1)-1:6*(NUM_NEIGHBOR_CELLS+1)];
assign enable_reading_2_4 = Local_enable_reading[8*(NUM_NEIGHBOR_CELLS+1)-1:7*(NUM_NEIGHBOR_CELLS+1)];
assign enable_reading_3_1 = Local_enable_reading[9*(NUM_NEIGHBOR_CELLS+1)-1:8*(NUM_NEIGHBOR_CELLS+1)];
assign enable_reading_3_2 = Local_enable_reading[10*(NUM_NEIGHBOR_CELLS+1)-1:9*(NUM_NEIGHBOR_CELLS+1)];
assign enable_reading_3_3 = Local_enable_reading[11*(NUM_NEIGHBOR_CELLS+1)-1:10*(NUM_NEIGHBOR_CELLS+1)];
assign enable_reading_3_4 = Local_enable_reading[12*(NUM_NEIGHBOR_CELLS+1)-1:11*(NUM_NEIGHBOR_CELLS+1)];
assign enable_reading_4_1 = Local_enable_reading[13*(NUM_NEIGHBOR_CELLS+1)-1:12*(NUM_NEIGHBOR_CELLS+1)];
assign enable_reading_4_2 = Local_enable_reading[14*(NUM_NEIGHBOR_CELLS+1)-1:13*(NUM_NEIGHBOR_CELLS+1)];
assign enable_reading_4_3 = Local_enable_reading[15*(NUM_NEIGHBOR_CELLS+1)-1:14*(NUM_NEIGHBOR_CELLS+1)];
assign enable_reading_4_4 = Local_enable_reading[16*(NUM_NEIGHBOR_CELLS+1)-1:15*(NUM_NEIGHBOR_CELLS+1)];

reg [NUM_NEIGHBOR_CELLS:0] reg_Cell_to_FSM_read_success_bit_1_1;
reg [NUM_NEIGHBOR_CELLS:0] reg_Cell_to_FSM_read_success_bit_1_2;
reg [NUM_NEIGHBOR_CELLS:0] reg_Cell_to_FSM_read_success_bit_1_3;
reg [NUM_NEIGHBOR_CELLS:0] reg_Cell_to_FSM_read_success_bit_1_4;
reg [NUM_NEIGHBOR_CELLS:0] reg_Cell_to_FSM_read_success_bit_2_1;
reg [NUM_NEIGHBOR_CELLS:0] reg_Cell_to_FSM_read_success_bit_2_2;
reg [NUM_NEIGHBOR_CELLS:0] reg_Cell_to_FSM_read_success_bit_2_3;
reg [NUM_NEIGHBOR_CELLS:0] reg_Cell_to_FSM_read_success_bit_2_4;
reg [NUM_NEIGHBOR_CELLS:0] reg_Cell_to_FSM_read_success_bit_3_1;
reg [NUM_NEIGHBOR_CELLS:0] reg_Cell_to_FSM_read_success_bit_3_2;
reg [NUM_NEIGHBOR_CELLS:0] reg_Cell_to_FSM_read_success_bit_3_3;
reg [NUM_NEIGHBOR_CELLS:0] reg_Cell_to_FSM_read_success_bit_3_4;
reg [NUM_NEIGHBOR_CELLS:0] reg_Cell_to_FSM_read_success_bit_4_1;
reg [NUM_NEIGHBOR_CELLS:0] reg_Cell_to_FSM_read_success_bit_4_2;
reg [NUM_NEIGHBOR_CELLS:0] reg_Cell_to_FSM_read_success_bit_4_3;
reg [NUM_NEIGHBOR_CELLS:0] reg_Cell_to_FSM_read_success_bit_4_4;
assign Cell_to_FSM_read_success_bit[1*(NUM_NEIGHBOR_CELLS+1)-1:0*(NUM_NEIGHBOR_CELLS+1)] = reg_Cell_to_FSM_read_success_bit_1_1;
assign Cell_to_FSM_read_success_bit[2*(NUM_NEIGHBOR_CELLS+1)-1:1*(NUM_NEIGHBOR_CELLS+1)] = reg_Cell_to_FSM_read_success_bit_1_2;
assign Cell_to_FSM_read_success_bit[3*(NUM_NEIGHBOR_CELLS+1)-1:2*(NUM_NEIGHBOR_CELLS+1)] = reg_Cell_to_FSM_read_success_bit_1_3;
assign Cell_to_FSM_read_success_bit[4*(NUM_NEIGHBOR_CELLS+1)-1:3*(NUM_NEIGHBOR_CELLS+1)] = reg_Cell_to_FSM_read_success_bit_1_4;
assign Cell_to_FSM_read_success_bit[5*(NUM_NEIGHBOR_CELLS+1)-1:4*(NUM_NEIGHBOR_CELLS+1)] = reg_Cell_to_FSM_read_success_bit_2_1;
assign Cell_to_FSM_read_success_bit[6*(NUM_NEIGHBOR_CELLS+1)-1:5*(NUM_NEIGHBOR_CELLS+1)] = reg_Cell_to_FSM_read_success_bit_2_2;
assign Cell_to_FSM_read_success_bit[7*(NUM_NEIGHBOR_CELLS+1)-1:6*(NUM_NEIGHBOR_CELLS+1)] = reg_Cell_to_FSM_read_success_bit_2_3;
assign Cell_to_FSM_read_success_bit[8*(NUM_NEIGHBOR_CELLS+1)-1:7*(NUM_NEIGHBOR_CELLS+1)] = reg_Cell_to_FSM_read_success_bit_2_4;
assign Cell_to_FSM_read_success_bit[9*(NUM_NEIGHBOR_CELLS+1)-1:8*(NUM_NEIGHBOR_CELLS+1)] = reg_Cell_to_FSM_read_success_bit_3_1;
assign Cell_to_FSM_read_success_bit[10*(NUM_NEIGHBOR_CELLS+1)-1:9*(NUM_NEIGHBOR_CELLS+1)] = reg_Cell_to_FSM_read_success_bit_3_2;
assign Cell_to_FSM_read_success_bit[11*(NUM_NEIGHBOR_CELLS+1)-1:10*(NUM_NEIGHBOR_CELLS+1)] = reg_Cell_to_FSM_read_success_bit_3_3;
assign Cell_to_FSM_read_success_bit[12*(NUM_NEIGHBOR_CELLS+1)-1:11*(NUM_NEIGHBOR_CELLS+1)] = reg_Cell_to_FSM_read_success_bit_3_4;
assign Cell_to_FSM_read_success_bit[13*(NUM_NEIGHBOR_CELLS+1)-1:12*(NUM_NEIGHBOR_CELLS+1)] = reg_Cell_to_FSM_read_success_bit_4_1;
assign Cell_to_FSM_read_success_bit[14*(NUM_NEIGHBOR_CELLS+1)-1:13*(NUM_NEIGHBOR_CELLS+1)] = reg_Cell_to_FSM_read_success_bit_4_2;
assign Cell_to_FSM_read_success_bit[15*(NUM_NEIGHBOR_CELLS+1)-1:14*(NUM_NEIGHBOR_CELLS+1)] = reg_Cell_to_FSM_read_success_bit_4_3;
assign Cell_to_FSM_read_success_bit[16*(NUM_NEIGHBOR_CELLS+1)-1:15*(NUM_NEIGHBOR_CELLS+1)] = reg_Cell_to_FSM_read_success_bit_4_4;

reg [TOTAL_CELL_NUM*CELL_ADDR_WIDTH-1:0] reg_FSM_to_Cell_read_addr;
assign FSM_to_Cell_read_addr = reg_FSM_to_Cell_read_addr;

wire [RDADDR_ARBITER_SIZE-1:0] arbiter_1_1_mid;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_1_2_mid;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_1_3_mid;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_1_4_mid;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_2_1_mid;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_2_2_mid;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_2_3_mid;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_2_4_mid;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_3_1_mid;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_3_2_mid;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_3_3_mid;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_3_4_mid;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_4_1_mid;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_4_2_mid;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_4_3_mid;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_4_4_mid;

wire [RDADDR_ARBITER_SIZE-1:0] arbiter_1_1_top;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_1_2_top;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_1_3_top;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_1_4_top;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_2_1_top;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_2_2_top;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_2_3_top;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_2_4_top;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_3_1_top;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_3_2_top;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_3_3_top;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_3_4_top;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_4_1_top;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_4_2_top;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_4_3_top;
wire [RDADDR_ARBITER_SIZE-1:0] arbiter_4_4_top;

wire [RDADDR_ARBITER_BOTTOM_SIZE-1:0] arbiter_1_1_bottom;
wire [RDADDR_ARBITER_BOTTOM_SIZE-1:0] arbiter_1_2_bottom;
wire [RDADDR_ARBITER_BOTTOM_SIZE-1:0] arbiter_1_3_bottom;
wire [RDADDR_ARBITER_BOTTOM_SIZE-1:0] arbiter_1_4_bottom;
wire [RDADDR_ARBITER_BOTTOM_SIZE-1:0] arbiter_2_1_bottom;
wire [RDADDR_ARBITER_BOTTOM_SIZE-1:0] arbiter_2_2_bottom;
wire [RDADDR_ARBITER_BOTTOM_SIZE-1:0] arbiter_2_3_bottom;
wire [RDADDR_ARBITER_BOTTOM_SIZE-1:0] arbiter_2_4_bottom;
wire [RDADDR_ARBITER_BOTTOM_SIZE-1:0] arbiter_3_1_bottom;
wire [RDADDR_ARBITER_BOTTOM_SIZE-1:0] arbiter_3_2_bottom;
wire [RDADDR_ARBITER_BOTTOM_SIZE-1:0] arbiter_3_3_bottom;
wire [RDADDR_ARBITER_BOTTOM_SIZE-1:0] arbiter_3_4_bottom;
wire [RDADDR_ARBITER_BOTTOM_SIZE-1:0] arbiter_4_1_bottom;
wire [RDADDR_ARBITER_BOTTOM_SIZE-1:0] arbiter_4_2_bottom;
wire [RDADDR_ARBITER_BOTTOM_SIZE-1:0] arbiter_4_3_bottom;
wire [RDADDR_ARBITER_BOTTOM_SIZE-1:0] arbiter_4_4_bottom;

always@(*)
	begin
	case (cellz)
		1: 
			begin
			if (arbiter_1_1_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_1_top[0])
				begin
				reg_FSM_to_Cell_read_addr[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_top[1])
				begin
				reg_FSM_to_Cell_read_addr[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_top[2])
				begin
				reg_FSM_to_Cell_read_addr[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_top[3])
				begin
				reg_FSM_to_Cell_read_addr[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_top[4])
				begin
				reg_FSM_to_Cell_read_addr[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH] = 0;
			if (arbiter_1_1_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_2_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_2_top[0])
				begin
				reg_FSM_to_Cell_read_addr[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_top[1])
				begin
				reg_FSM_to_Cell_read_addr[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_top[2])
				begin
				reg_FSM_to_Cell_read_addr[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_top[3])
				begin
				reg_FSM_to_Cell_read_addr[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_top[4])
				begin
				reg_FSM_to_Cell_read_addr[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH] = 0;
			if (arbiter_1_2_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_3_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_3_top[0])
				begin
				reg_FSM_to_Cell_read_addr[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_top[1])
				begin
				reg_FSM_to_Cell_read_addr[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_top[2])
				begin
				reg_FSM_to_Cell_read_addr[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_top[3])
				begin
				reg_FSM_to_Cell_read_addr[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_top[4])
				begin
				reg_FSM_to_Cell_read_addr[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH] = 0;
			if (arbiter_1_3_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_4_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_4_top[0])
				begin
				reg_FSM_to_Cell_read_addr[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_top[1])
				begin
				reg_FSM_to_Cell_read_addr[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_top[2])
				begin
				reg_FSM_to_Cell_read_addr[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_top[3])
				begin
				reg_FSM_to_Cell_read_addr[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_top[4])
				begin
				reg_FSM_to_Cell_read_addr[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[15*CELL_ADDR_WIDTH-1:14*CELL_ADDR_WIDTH] = 0;
			if (arbiter_1_4_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[16*CELL_ADDR_WIDTH-1:15*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[16*CELL_ADDR_WIDTH-1:15*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[16*CELL_ADDR_WIDTH-1:15*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[16*CELL_ADDR_WIDTH-1:15*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[16*CELL_ADDR_WIDTH-1:15*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_1_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[17*CELL_ADDR_WIDTH-1:16*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[17*CELL_ADDR_WIDTH-1:16*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[17*CELL_ADDR_WIDTH-1:16*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[17*CELL_ADDR_WIDTH-1:16*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[17*CELL_ADDR_WIDTH-1:16*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[17*CELL_ADDR_WIDTH-1:16*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_1_top[0])
				begin
				reg_FSM_to_Cell_read_addr[18*CELL_ADDR_WIDTH-1:17*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_top[1])
				begin
				reg_FSM_to_Cell_read_addr[18*CELL_ADDR_WIDTH-1:17*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_top[2])
				begin
				reg_FSM_to_Cell_read_addr[18*CELL_ADDR_WIDTH-1:17*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_top[3])
				begin
				reg_FSM_to_Cell_read_addr[18*CELL_ADDR_WIDTH-1:17*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_top[4])
				begin
				reg_FSM_to_Cell_read_addr[18*CELL_ADDR_WIDTH-1:17*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[18*CELL_ADDR_WIDTH-1:17*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[19*CELL_ADDR_WIDTH-1:18*CELL_ADDR_WIDTH] = 0;
			if (arbiter_2_1_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[20*CELL_ADDR_WIDTH-1:19*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[20*CELL_ADDR_WIDTH-1:19*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[20*CELL_ADDR_WIDTH-1:19*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[20*CELL_ADDR_WIDTH-1:19*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[20*CELL_ADDR_WIDTH-1:19*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_2_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[21*CELL_ADDR_WIDTH-1:20*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[21*CELL_ADDR_WIDTH-1:20*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[21*CELL_ADDR_WIDTH-1:20*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[21*CELL_ADDR_WIDTH-1:20*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[21*CELL_ADDR_WIDTH-1:20*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[21*CELL_ADDR_WIDTH-1:20*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_2_top[0])
				begin
				reg_FSM_to_Cell_read_addr[22*CELL_ADDR_WIDTH-1:21*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_top[1])
				begin
				reg_FSM_to_Cell_read_addr[22*CELL_ADDR_WIDTH-1:21*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_top[2])
				begin
				reg_FSM_to_Cell_read_addr[22*CELL_ADDR_WIDTH-1:21*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_top[3])
				begin
				reg_FSM_to_Cell_read_addr[22*CELL_ADDR_WIDTH-1:21*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_top[4])
				begin
				reg_FSM_to_Cell_read_addr[22*CELL_ADDR_WIDTH-1:21*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[22*CELL_ADDR_WIDTH-1:21*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[23*CELL_ADDR_WIDTH-1:22*CELL_ADDR_WIDTH] = 0;
			if (arbiter_2_2_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[24*CELL_ADDR_WIDTH-1:23*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[24*CELL_ADDR_WIDTH-1:23*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[24*CELL_ADDR_WIDTH-1:23*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[24*CELL_ADDR_WIDTH-1:23*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[24*CELL_ADDR_WIDTH-1:23*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_3_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[25*CELL_ADDR_WIDTH-1:24*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[25*CELL_ADDR_WIDTH-1:24*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[25*CELL_ADDR_WIDTH-1:24*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[25*CELL_ADDR_WIDTH-1:24*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[25*CELL_ADDR_WIDTH-1:24*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[25*CELL_ADDR_WIDTH-1:24*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_3_top[0])
				begin
				reg_FSM_to_Cell_read_addr[26*CELL_ADDR_WIDTH-1:25*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_top[1])
				begin
				reg_FSM_to_Cell_read_addr[26*CELL_ADDR_WIDTH-1:25*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_top[2])
				begin
				reg_FSM_to_Cell_read_addr[26*CELL_ADDR_WIDTH-1:25*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_top[3])
				begin
				reg_FSM_to_Cell_read_addr[26*CELL_ADDR_WIDTH-1:25*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_top[4])
				begin
				reg_FSM_to_Cell_read_addr[26*CELL_ADDR_WIDTH-1:25*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[26*CELL_ADDR_WIDTH-1:25*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[27*CELL_ADDR_WIDTH-1:26*CELL_ADDR_WIDTH] = 0;
			if (arbiter_2_3_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[28*CELL_ADDR_WIDTH-1:27*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[28*CELL_ADDR_WIDTH-1:27*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[28*CELL_ADDR_WIDTH-1:27*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[28*CELL_ADDR_WIDTH-1:27*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[28*CELL_ADDR_WIDTH-1:27*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_4_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[29*CELL_ADDR_WIDTH-1:28*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[29*CELL_ADDR_WIDTH-1:28*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[29*CELL_ADDR_WIDTH-1:28*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[29*CELL_ADDR_WIDTH-1:28*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[29*CELL_ADDR_WIDTH-1:28*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[29*CELL_ADDR_WIDTH-1:28*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_4_top[0])
				begin
				reg_FSM_to_Cell_read_addr[30*CELL_ADDR_WIDTH-1:29*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_top[1])
				begin
				reg_FSM_to_Cell_read_addr[30*CELL_ADDR_WIDTH-1:29*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_top[2])
				begin
				reg_FSM_to_Cell_read_addr[30*CELL_ADDR_WIDTH-1:29*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_top[3])
				begin
				reg_FSM_to_Cell_read_addr[30*CELL_ADDR_WIDTH-1:29*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_top[4])
				begin
				reg_FSM_to_Cell_read_addr[30*CELL_ADDR_WIDTH-1:29*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[30*CELL_ADDR_WIDTH-1:29*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[31*CELL_ADDR_WIDTH-1:30*CELL_ADDR_WIDTH] = 0;
			if (arbiter_2_4_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[32*CELL_ADDR_WIDTH-1:31*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[32*CELL_ADDR_WIDTH-1:31*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[32*CELL_ADDR_WIDTH-1:31*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[32*CELL_ADDR_WIDTH-1:31*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[32*CELL_ADDR_WIDTH-1:31*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_1_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[33*CELL_ADDR_WIDTH-1:32*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[33*CELL_ADDR_WIDTH-1:32*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[33*CELL_ADDR_WIDTH-1:32*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[33*CELL_ADDR_WIDTH-1:32*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[33*CELL_ADDR_WIDTH-1:32*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[33*CELL_ADDR_WIDTH-1:32*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_1_top[0])
				begin
				reg_FSM_to_Cell_read_addr[34*CELL_ADDR_WIDTH-1:33*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_top[1])
				begin
				reg_FSM_to_Cell_read_addr[34*CELL_ADDR_WIDTH-1:33*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_top[2])
				begin
				reg_FSM_to_Cell_read_addr[34*CELL_ADDR_WIDTH-1:33*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_top[3])
				begin
				reg_FSM_to_Cell_read_addr[34*CELL_ADDR_WIDTH-1:33*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_top[4])
				begin
				reg_FSM_to_Cell_read_addr[34*CELL_ADDR_WIDTH-1:33*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[34*CELL_ADDR_WIDTH-1:33*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[35*CELL_ADDR_WIDTH-1:34*CELL_ADDR_WIDTH] = 0;
			if (arbiter_3_1_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[36*CELL_ADDR_WIDTH-1:35*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[36*CELL_ADDR_WIDTH-1:35*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[36*CELL_ADDR_WIDTH-1:35*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[36*CELL_ADDR_WIDTH-1:35*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[36*CELL_ADDR_WIDTH-1:35*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_2_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[37*CELL_ADDR_WIDTH-1:36*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[37*CELL_ADDR_WIDTH-1:36*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[37*CELL_ADDR_WIDTH-1:36*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[37*CELL_ADDR_WIDTH-1:36*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[37*CELL_ADDR_WIDTH-1:36*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[37*CELL_ADDR_WIDTH-1:36*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_2_top[0])
				begin
				reg_FSM_to_Cell_read_addr[38*CELL_ADDR_WIDTH-1:37*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_top[1])
				begin
				reg_FSM_to_Cell_read_addr[38*CELL_ADDR_WIDTH-1:37*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_top[2])
				begin
				reg_FSM_to_Cell_read_addr[38*CELL_ADDR_WIDTH-1:37*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_top[3])
				begin
				reg_FSM_to_Cell_read_addr[38*CELL_ADDR_WIDTH-1:37*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_top[4])
				begin
				reg_FSM_to_Cell_read_addr[38*CELL_ADDR_WIDTH-1:37*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[38*CELL_ADDR_WIDTH-1:37*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[39*CELL_ADDR_WIDTH-1:38*CELL_ADDR_WIDTH] = 0;
			if (arbiter_3_2_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[40*CELL_ADDR_WIDTH-1:39*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[40*CELL_ADDR_WIDTH-1:39*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[40*CELL_ADDR_WIDTH-1:39*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[40*CELL_ADDR_WIDTH-1:39*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[40*CELL_ADDR_WIDTH-1:39*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_3_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[41*CELL_ADDR_WIDTH-1:40*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[41*CELL_ADDR_WIDTH-1:40*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[41*CELL_ADDR_WIDTH-1:40*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[41*CELL_ADDR_WIDTH-1:40*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[41*CELL_ADDR_WIDTH-1:40*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[41*CELL_ADDR_WIDTH-1:40*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_3_top[0])
				begin
				reg_FSM_to_Cell_read_addr[42*CELL_ADDR_WIDTH-1:41*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_top[1])
				begin
				reg_FSM_to_Cell_read_addr[42*CELL_ADDR_WIDTH-1:41*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_top[2])
				begin
				reg_FSM_to_Cell_read_addr[42*CELL_ADDR_WIDTH-1:41*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_top[3])
				begin
				reg_FSM_to_Cell_read_addr[42*CELL_ADDR_WIDTH-1:41*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_top[4])
				begin
				reg_FSM_to_Cell_read_addr[42*CELL_ADDR_WIDTH-1:41*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[42*CELL_ADDR_WIDTH-1:41*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[43*CELL_ADDR_WIDTH-1:42*CELL_ADDR_WIDTH] = 0;
			if (arbiter_3_3_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[44*CELL_ADDR_WIDTH-1:43*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[44*CELL_ADDR_WIDTH-1:43*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[44*CELL_ADDR_WIDTH-1:43*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[44*CELL_ADDR_WIDTH-1:43*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[44*CELL_ADDR_WIDTH-1:43*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_4_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[45*CELL_ADDR_WIDTH-1:44*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[45*CELL_ADDR_WIDTH-1:44*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[45*CELL_ADDR_WIDTH-1:44*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[45*CELL_ADDR_WIDTH-1:44*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[45*CELL_ADDR_WIDTH-1:44*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[45*CELL_ADDR_WIDTH-1:44*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_4_top[0])
				begin
				reg_FSM_to_Cell_read_addr[46*CELL_ADDR_WIDTH-1:45*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_top[1])
				begin
				reg_FSM_to_Cell_read_addr[46*CELL_ADDR_WIDTH-1:45*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_top[2])
				begin
				reg_FSM_to_Cell_read_addr[46*CELL_ADDR_WIDTH-1:45*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_top[3])
				begin
				reg_FSM_to_Cell_read_addr[46*CELL_ADDR_WIDTH-1:45*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_top[4])
				begin
				reg_FSM_to_Cell_read_addr[46*CELL_ADDR_WIDTH-1:45*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[46*CELL_ADDR_WIDTH-1:45*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[47*CELL_ADDR_WIDTH-1:46*CELL_ADDR_WIDTH] = 0;
			if (arbiter_3_4_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[48*CELL_ADDR_WIDTH-1:47*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[48*CELL_ADDR_WIDTH-1:47*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[48*CELL_ADDR_WIDTH-1:47*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[48*CELL_ADDR_WIDTH-1:47*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[48*CELL_ADDR_WIDTH-1:47*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_1_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[49*CELL_ADDR_WIDTH-1:48*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[49*CELL_ADDR_WIDTH-1:48*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[49*CELL_ADDR_WIDTH-1:48*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[49*CELL_ADDR_WIDTH-1:48*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[49*CELL_ADDR_WIDTH-1:48*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[49*CELL_ADDR_WIDTH-1:48*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_1_top[0])
				begin
				reg_FSM_to_Cell_read_addr[50*CELL_ADDR_WIDTH-1:49*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_top[1])
				begin
				reg_FSM_to_Cell_read_addr[50*CELL_ADDR_WIDTH-1:49*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_top[2])
				begin
				reg_FSM_to_Cell_read_addr[50*CELL_ADDR_WIDTH-1:49*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_top[3])
				begin
				reg_FSM_to_Cell_read_addr[50*CELL_ADDR_WIDTH-1:49*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_top[4])
				begin
				reg_FSM_to_Cell_read_addr[50*CELL_ADDR_WIDTH-1:49*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[50*CELL_ADDR_WIDTH-1:49*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[51*CELL_ADDR_WIDTH-1:50*CELL_ADDR_WIDTH] = 0;
			if (arbiter_4_1_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[52*CELL_ADDR_WIDTH-1:51*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[52*CELL_ADDR_WIDTH-1:51*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[52*CELL_ADDR_WIDTH-1:51*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[52*CELL_ADDR_WIDTH-1:51*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[52*CELL_ADDR_WIDTH-1:51*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_2_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[53*CELL_ADDR_WIDTH-1:52*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[53*CELL_ADDR_WIDTH-1:52*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[53*CELL_ADDR_WIDTH-1:52*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[53*CELL_ADDR_WIDTH-1:52*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[53*CELL_ADDR_WIDTH-1:52*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[53*CELL_ADDR_WIDTH-1:52*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_2_top[0])
				begin
				reg_FSM_to_Cell_read_addr[54*CELL_ADDR_WIDTH-1:53*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_top[1])
				begin
				reg_FSM_to_Cell_read_addr[54*CELL_ADDR_WIDTH-1:53*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_top[2])
				begin
				reg_FSM_to_Cell_read_addr[54*CELL_ADDR_WIDTH-1:53*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_top[3])
				begin
				reg_FSM_to_Cell_read_addr[54*CELL_ADDR_WIDTH-1:53*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_top[4])
				begin
				reg_FSM_to_Cell_read_addr[54*CELL_ADDR_WIDTH-1:53*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[54*CELL_ADDR_WIDTH-1:53*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[55*CELL_ADDR_WIDTH-1:54*CELL_ADDR_WIDTH] = 0;
			if (arbiter_4_2_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[56*CELL_ADDR_WIDTH-1:55*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[56*CELL_ADDR_WIDTH-1:55*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[56*CELL_ADDR_WIDTH-1:55*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[56*CELL_ADDR_WIDTH-1:55*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[56*CELL_ADDR_WIDTH-1:55*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_3_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[57*CELL_ADDR_WIDTH-1:56*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[57*CELL_ADDR_WIDTH-1:56*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[57*CELL_ADDR_WIDTH-1:56*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[57*CELL_ADDR_WIDTH-1:56*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[57*CELL_ADDR_WIDTH-1:56*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[57*CELL_ADDR_WIDTH-1:56*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_3_top[0])
				begin
				reg_FSM_to_Cell_read_addr[58*CELL_ADDR_WIDTH-1:57*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_top[1])
				begin
				reg_FSM_to_Cell_read_addr[58*CELL_ADDR_WIDTH-1:57*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_top[2])
				begin
				reg_FSM_to_Cell_read_addr[58*CELL_ADDR_WIDTH-1:57*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_top[3])
				begin
				reg_FSM_to_Cell_read_addr[58*CELL_ADDR_WIDTH-1:57*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_top[4])
				begin
				reg_FSM_to_Cell_read_addr[58*CELL_ADDR_WIDTH-1:57*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[58*CELL_ADDR_WIDTH-1:57*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[59*CELL_ADDR_WIDTH-1:58*CELL_ADDR_WIDTH] = 0;
			if (arbiter_4_3_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[60*CELL_ADDR_WIDTH-1:59*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[60*CELL_ADDR_WIDTH-1:59*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[60*CELL_ADDR_WIDTH-1:59*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[60*CELL_ADDR_WIDTH-1:59*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[60*CELL_ADDR_WIDTH-1:59*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_4_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[61*CELL_ADDR_WIDTH-1:60*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[61*CELL_ADDR_WIDTH-1:60*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[61*CELL_ADDR_WIDTH-1:60*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[61*CELL_ADDR_WIDTH-1:60*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[61*CELL_ADDR_WIDTH-1:60*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[61*CELL_ADDR_WIDTH-1:60*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_4_top[0])
				begin
				reg_FSM_to_Cell_read_addr[62*CELL_ADDR_WIDTH-1:61*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_top[1])
				begin
				reg_FSM_to_Cell_read_addr[62*CELL_ADDR_WIDTH-1:61*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_top[2])
				begin
				reg_FSM_to_Cell_read_addr[62*CELL_ADDR_WIDTH-1:61*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_top[3])
				begin
				reg_FSM_to_Cell_read_addr[62*CELL_ADDR_WIDTH-1:61*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_top[4])
				begin
				reg_FSM_to_Cell_read_addr[62*CELL_ADDR_WIDTH-1:61*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[62*CELL_ADDR_WIDTH-1:61*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[63*CELL_ADDR_WIDTH-1:62*CELL_ADDR_WIDTH] = 0;
			if (arbiter_4_4_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[64*CELL_ADDR_WIDTH-1:63*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[64*CELL_ADDR_WIDTH-1:63*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[64*CELL_ADDR_WIDTH-1:63*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[64*CELL_ADDR_WIDTH-1:63*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[64*CELL_ADDR_WIDTH-1:63*CELL_ADDR_WIDTH] = 0;
				end
			end
		2:
			begin
			if (arbiter_1_1_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_1_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_1_top[0])
				begin
				reg_FSM_to_Cell_read_addr[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_top[1])
				begin
				reg_FSM_to_Cell_read_addr[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_top[2])
				begin
				reg_FSM_to_Cell_read_addr[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_top[3])
				begin
				reg_FSM_to_Cell_read_addr[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_top[4])
				begin
				reg_FSM_to_Cell_read_addr[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH] = 0;
			if (arbiter_1_2_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_2_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_2_top[0])
				begin
				reg_FSM_to_Cell_read_addr[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_top[1])
				begin
				reg_FSM_to_Cell_read_addr[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_top[2])
				begin
				reg_FSM_to_Cell_read_addr[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_top[3])
				begin
				reg_FSM_to_Cell_read_addr[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_top[4])
				begin
				reg_FSM_to_Cell_read_addr[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH] = 0;
			if (arbiter_1_3_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_3_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_3_top[0])
				begin
				reg_FSM_to_Cell_read_addr[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_top[1])
				begin
				reg_FSM_to_Cell_read_addr[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_top[2])
				begin
				reg_FSM_to_Cell_read_addr[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_top[3])
				begin
				reg_FSM_to_Cell_read_addr[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_top[4])
				begin
				reg_FSM_to_Cell_read_addr[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH] = 0;
			if (arbiter_1_4_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_4_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_4_top[0])
				begin
				reg_FSM_to_Cell_read_addr[15*CELL_ADDR_WIDTH-1:14*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_top[1])
				begin
				reg_FSM_to_Cell_read_addr[15*CELL_ADDR_WIDTH-1:14*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_top[2])
				begin
				reg_FSM_to_Cell_read_addr[15*CELL_ADDR_WIDTH-1:14*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_top[3])
				begin
				reg_FSM_to_Cell_read_addr[15*CELL_ADDR_WIDTH-1:14*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_top[4])
				begin
				reg_FSM_to_Cell_read_addr[15*CELL_ADDR_WIDTH-1:14*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[15*CELL_ADDR_WIDTH-1:14*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[16*CELL_ADDR_WIDTH-1:15*CELL_ADDR_WIDTH] = 0;
			if (arbiter_2_1_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[17*CELL_ADDR_WIDTH-1:16*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[17*CELL_ADDR_WIDTH-1:16*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[17*CELL_ADDR_WIDTH-1:16*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[17*CELL_ADDR_WIDTH-1:16*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[17*CELL_ADDR_WIDTH-1:16*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_1_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[18*CELL_ADDR_WIDTH-1:17*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[18*CELL_ADDR_WIDTH-1:17*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[18*CELL_ADDR_WIDTH-1:17*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[18*CELL_ADDR_WIDTH-1:17*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[18*CELL_ADDR_WIDTH-1:17*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[18*CELL_ADDR_WIDTH-1:17*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_1_top[0])
				begin
				reg_FSM_to_Cell_read_addr[19*CELL_ADDR_WIDTH-1:18*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_top[1])
				begin
				reg_FSM_to_Cell_read_addr[19*CELL_ADDR_WIDTH-1:18*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_top[2])
				begin
				reg_FSM_to_Cell_read_addr[19*CELL_ADDR_WIDTH-1:18*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_top[3])
				begin
				reg_FSM_to_Cell_read_addr[19*CELL_ADDR_WIDTH-1:18*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_top[4])
				begin
				reg_FSM_to_Cell_read_addr[19*CELL_ADDR_WIDTH-1:18*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[19*CELL_ADDR_WIDTH-1:18*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[20*CELL_ADDR_WIDTH-1:19*CELL_ADDR_WIDTH] = 0;
			if (arbiter_2_2_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[21*CELL_ADDR_WIDTH-1:20*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[21*CELL_ADDR_WIDTH-1:20*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[21*CELL_ADDR_WIDTH-1:20*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[21*CELL_ADDR_WIDTH-1:20*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[21*CELL_ADDR_WIDTH-1:20*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_2_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[22*CELL_ADDR_WIDTH-1:21*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[22*CELL_ADDR_WIDTH-1:21*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[22*CELL_ADDR_WIDTH-1:21*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[22*CELL_ADDR_WIDTH-1:21*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[22*CELL_ADDR_WIDTH-1:21*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[22*CELL_ADDR_WIDTH-1:21*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_2_top[0])
				begin
				reg_FSM_to_Cell_read_addr[23*CELL_ADDR_WIDTH-1:22*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_top[1])
				begin
				reg_FSM_to_Cell_read_addr[23*CELL_ADDR_WIDTH-1:22*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_top[2])
				begin
				reg_FSM_to_Cell_read_addr[23*CELL_ADDR_WIDTH-1:22*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_top[3])
				begin
				reg_FSM_to_Cell_read_addr[23*CELL_ADDR_WIDTH-1:22*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_top[4])
				begin
				reg_FSM_to_Cell_read_addr[23*CELL_ADDR_WIDTH-1:22*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[23*CELL_ADDR_WIDTH-1:22*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[24*CELL_ADDR_WIDTH-1:23*CELL_ADDR_WIDTH] = 0;
			if (arbiter_2_3_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[25*CELL_ADDR_WIDTH-1:24*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[25*CELL_ADDR_WIDTH-1:24*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[25*CELL_ADDR_WIDTH-1:24*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[25*CELL_ADDR_WIDTH-1:24*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[25*CELL_ADDR_WIDTH-1:24*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_3_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[26*CELL_ADDR_WIDTH-1:25*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[26*CELL_ADDR_WIDTH-1:25*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[26*CELL_ADDR_WIDTH-1:25*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[26*CELL_ADDR_WIDTH-1:25*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[26*CELL_ADDR_WIDTH-1:25*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[26*CELL_ADDR_WIDTH-1:25*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_3_top[0])
				begin
				reg_FSM_to_Cell_read_addr[27*CELL_ADDR_WIDTH-1:26*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_top[1])
				begin
				reg_FSM_to_Cell_read_addr[27*CELL_ADDR_WIDTH-1:26*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_top[2])
				begin
				reg_FSM_to_Cell_read_addr[27*CELL_ADDR_WIDTH-1:26*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_top[3])
				begin
				reg_FSM_to_Cell_read_addr[27*CELL_ADDR_WIDTH-1:26*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_top[4])
				begin
				reg_FSM_to_Cell_read_addr[27*CELL_ADDR_WIDTH-1:26*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[27*CELL_ADDR_WIDTH-1:26*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[28*CELL_ADDR_WIDTH-1:27*CELL_ADDR_WIDTH] = 0;
			if (arbiter_2_4_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[29*CELL_ADDR_WIDTH-1:28*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[29*CELL_ADDR_WIDTH-1:28*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[29*CELL_ADDR_WIDTH-1:28*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[29*CELL_ADDR_WIDTH-1:28*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[29*CELL_ADDR_WIDTH-1:28*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_4_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[30*CELL_ADDR_WIDTH-1:29*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[30*CELL_ADDR_WIDTH-1:29*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[30*CELL_ADDR_WIDTH-1:29*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[30*CELL_ADDR_WIDTH-1:29*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[30*CELL_ADDR_WIDTH-1:29*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[30*CELL_ADDR_WIDTH-1:29*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_4_top[0])
				begin
				reg_FSM_to_Cell_read_addr[31*CELL_ADDR_WIDTH-1:30*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_top[1])
				begin
				reg_FSM_to_Cell_read_addr[31*CELL_ADDR_WIDTH-1:30*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_top[2])
				begin
				reg_FSM_to_Cell_read_addr[31*CELL_ADDR_WIDTH-1:30*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_top[3])
				begin
				reg_FSM_to_Cell_read_addr[31*CELL_ADDR_WIDTH-1:30*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_top[4])
				begin
				reg_FSM_to_Cell_read_addr[31*CELL_ADDR_WIDTH-1:30*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[31*CELL_ADDR_WIDTH-1:30*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[32*CELL_ADDR_WIDTH-1:31*CELL_ADDR_WIDTH] = 0;
			if (arbiter_3_1_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[33*CELL_ADDR_WIDTH-1:32*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[33*CELL_ADDR_WIDTH-1:32*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[33*CELL_ADDR_WIDTH-1:32*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[33*CELL_ADDR_WIDTH-1:32*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[33*CELL_ADDR_WIDTH-1:32*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_1_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[34*CELL_ADDR_WIDTH-1:33*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[34*CELL_ADDR_WIDTH-1:33*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[34*CELL_ADDR_WIDTH-1:33*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[34*CELL_ADDR_WIDTH-1:33*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[34*CELL_ADDR_WIDTH-1:33*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[34*CELL_ADDR_WIDTH-1:33*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_1_top[0])
				begin
				reg_FSM_to_Cell_read_addr[35*CELL_ADDR_WIDTH-1:34*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_top[1])
				begin
				reg_FSM_to_Cell_read_addr[35*CELL_ADDR_WIDTH-1:34*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_top[2])
				begin
				reg_FSM_to_Cell_read_addr[35*CELL_ADDR_WIDTH-1:34*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_top[3])
				begin
				reg_FSM_to_Cell_read_addr[35*CELL_ADDR_WIDTH-1:34*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_top[4])
				begin
				reg_FSM_to_Cell_read_addr[35*CELL_ADDR_WIDTH-1:34*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[35*CELL_ADDR_WIDTH-1:34*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[36*CELL_ADDR_WIDTH-1:35*CELL_ADDR_WIDTH] = 0;
			if (arbiter_3_2_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[37*CELL_ADDR_WIDTH-1:36*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[37*CELL_ADDR_WIDTH-1:36*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[37*CELL_ADDR_WIDTH-1:36*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[37*CELL_ADDR_WIDTH-1:36*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[37*CELL_ADDR_WIDTH-1:36*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_2_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[38*CELL_ADDR_WIDTH-1:37*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[38*CELL_ADDR_WIDTH-1:37*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[38*CELL_ADDR_WIDTH-1:37*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[38*CELL_ADDR_WIDTH-1:37*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[38*CELL_ADDR_WIDTH-1:37*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[38*CELL_ADDR_WIDTH-1:37*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_2_top[0])
				begin
				reg_FSM_to_Cell_read_addr[39*CELL_ADDR_WIDTH-1:38*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_top[1])
				begin
				reg_FSM_to_Cell_read_addr[39*CELL_ADDR_WIDTH-1:38*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_top[2])
				begin
				reg_FSM_to_Cell_read_addr[39*CELL_ADDR_WIDTH-1:38*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_top[3])
				begin
				reg_FSM_to_Cell_read_addr[39*CELL_ADDR_WIDTH-1:38*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_top[4])
				begin
				reg_FSM_to_Cell_read_addr[39*CELL_ADDR_WIDTH-1:38*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[39*CELL_ADDR_WIDTH-1:38*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[40*CELL_ADDR_WIDTH-1:39*CELL_ADDR_WIDTH] = 0;
			if (arbiter_3_3_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[41*CELL_ADDR_WIDTH-1:40*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[41*CELL_ADDR_WIDTH-1:40*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[41*CELL_ADDR_WIDTH-1:40*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[41*CELL_ADDR_WIDTH-1:40*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[41*CELL_ADDR_WIDTH-1:40*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_3_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[42*CELL_ADDR_WIDTH-1:41*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[42*CELL_ADDR_WIDTH-1:41*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[42*CELL_ADDR_WIDTH-1:41*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[42*CELL_ADDR_WIDTH-1:41*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[42*CELL_ADDR_WIDTH-1:41*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[42*CELL_ADDR_WIDTH-1:41*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_3_top[0])
				begin
				reg_FSM_to_Cell_read_addr[43*CELL_ADDR_WIDTH-1:42*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_top[1])
				begin
				reg_FSM_to_Cell_read_addr[43*CELL_ADDR_WIDTH-1:42*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_top[2])
				begin
				reg_FSM_to_Cell_read_addr[43*CELL_ADDR_WIDTH-1:42*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_top[3])
				begin
				reg_FSM_to_Cell_read_addr[43*CELL_ADDR_WIDTH-1:42*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_top[4])
				begin
				reg_FSM_to_Cell_read_addr[43*CELL_ADDR_WIDTH-1:42*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[43*CELL_ADDR_WIDTH-1:42*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[44*CELL_ADDR_WIDTH-1:43*CELL_ADDR_WIDTH] = 0;
			if (arbiter_3_4_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[45*CELL_ADDR_WIDTH-1:44*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[45*CELL_ADDR_WIDTH-1:44*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[45*CELL_ADDR_WIDTH-1:44*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[45*CELL_ADDR_WIDTH-1:44*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[45*CELL_ADDR_WIDTH-1:44*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_4_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[46*CELL_ADDR_WIDTH-1:45*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[46*CELL_ADDR_WIDTH-1:45*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[46*CELL_ADDR_WIDTH-1:45*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[46*CELL_ADDR_WIDTH-1:45*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[46*CELL_ADDR_WIDTH-1:45*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[46*CELL_ADDR_WIDTH-1:45*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_4_top[0])
				begin
				reg_FSM_to_Cell_read_addr[47*CELL_ADDR_WIDTH-1:46*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_top[1])
				begin
				reg_FSM_to_Cell_read_addr[47*CELL_ADDR_WIDTH-1:46*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_top[2])
				begin
				reg_FSM_to_Cell_read_addr[47*CELL_ADDR_WIDTH-1:46*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_top[3])
				begin
				reg_FSM_to_Cell_read_addr[47*CELL_ADDR_WIDTH-1:46*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_top[4])
				begin
				reg_FSM_to_Cell_read_addr[47*CELL_ADDR_WIDTH-1:46*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[47*CELL_ADDR_WIDTH-1:46*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[48*CELL_ADDR_WIDTH-1:47*CELL_ADDR_WIDTH] = 0;
			if (arbiter_4_1_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[49*CELL_ADDR_WIDTH-1:48*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[49*CELL_ADDR_WIDTH-1:48*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[49*CELL_ADDR_WIDTH-1:48*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[49*CELL_ADDR_WIDTH-1:48*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[49*CELL_ADDR_WIDTH-1:48*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_1_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[50*CELL_ADDR_WIDTH-1:49*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[50*CELL_ADDR_WIDTH-1:49*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[50*CELL_ADDR_WIDTH-1:49*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[50*CELL_ADDR_WIDTH-1:49*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[50*CELL_ADDR_WIDTH-1:49*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[50*CELL_ADDR_WIDTH-1:49*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_1_top[0])
				begin
				reg_FSM_to_Cell_read_addr[51*CELL_ADDR_WIDTH-1:50*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_top[1])
				begin
				reg_FSM_to_Cell_read_addr[51*CELL_ADDR_WIDTH-1:50*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_top[2])
				begin
				reg_FSM_to_Cell_read_addr[51*CELL_ADDR_WIDTH-1:50*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_top[3])
				begin
				reg_FSM_to_Cell_read_addr[51*CELL_ADDR_WIDTH-1:50*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_top[4])
				begin
				reg_FSM_to_Cell_read_addr[51*CELL_ADDR_WIDTH-1:50*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[51*CELL_ADDR_WIDTH-1:50*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[52*CELL_ADDR_WIDTH-1:51*CELL_ADDR_WIDTH] = 0;
			if (arbiter_4_2_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[53*CELL_ADDR_WIDTH-1:52*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[53*CELL_ADDR_WIDTH-1:52*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[53*CELL_ADDR_WIDTH-1:52*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[53*CELL_ADDR_WIDTH-1:52*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[53*CELL_ADDR_WIDTH-1:52*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_2_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[54*CELL_ADDR_WIDTH-1:53*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[54*CELL_ADDR_WIDTH-1:53*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[54*CELL_ADDR_WIDTH-1:53*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[54*CELL_ADDR_WIDTH-1:53*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[54*CELL_ADDR_WIDTH-1:53*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[54*CELL_ADDR_WIDTH-1:53*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_2_top[0])
				begin
				reg_FSM_to_Cell_read_addr[55*CELL_ADDR_WIDTH-1:54*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_top[1])
				begin
				reg_FSM_to_Cell_read_addr[55*CELL_ADDR_WIDTH-1:54*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_top[2])
				begin
				reg_FSM_to_Cell_read_addr[55*CELL_ADDR_WIDTH-1:54*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_top[3])
				begin
				reg_FSM_to_Cell_read_addr[55*CELL_ADDR_WIDTH-1:54*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_top[4])
				begin
				reg_FSM_to_Cell_read_addr[55*CELL_ADDR_WIDTH-1:54*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[55*CELL_ADDR_WIDTH-1:54*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[56*CELL_ADDR_WIDTH-1:55*CELL_ADDR_WIDTH] = 0;
			if (arbiter_4_3_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[57*CELL_ADDR_WIDTH-1:56*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[57*CELL_ADDR_WIDTH-1:56*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[57*CELL_ADDR_WIDTH-1:56*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[57*CELL_ADDR_WIDTH-1:56*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[57*CELL_ADDR_WIDTH-1:56*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_3_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[58*CELL_ADDR_WIDTH-1:57*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[58*CELL_ADDR_WIDTH-1:57*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[58*CELL_ADDR_WIDTH-1:57*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[58*CELL_ADDR_WIDTH-1:57*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[58*CELL_ADDR_WIDTH-1:57*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[58*CELL_ADDR_WIDTH-1:57*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_3_top[0])
				begin
				reg_FSM_to_Cell_read_addr[59*CELL_ADDR_WIDTH-1:58*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_top[1])
				begin
				reg_FSM_to_Cell_read_addr[59*CELL_ADDR_WIDTH-1:58*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_top[2])
				begin
				reg_FSM_to_Cell_read_addr[59*CELL_ADDR_WIDTH-1:58*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_top[3])
				begin
				reg_FSM_to_Cell_read_addr[59*CELL_ADDR_WIDTH-1:58*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_top[4])
				begin
				reg_FSM_to_Cell_read_addr[59*CELL_ADDR_WIDTH-1:58*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[59*CELL_ADDR_WIDTH-1:58*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[60*CELL_ADDR_WIDTH-1:59*CELL_ADDR_WIDTH] = 0;
			if (arbiter_4_4_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[61*CELL_ADDR_WIDTH-1:60*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[61*CELL_ADDR_WIDTH-1:60*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[61*CELL_ADDR_WIDTH-1:60*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[61*CELL_ADDR_WIDTH-1:60*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[61*CELL_ADDR_WIDTH-1:60*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_4_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[62*CELL_ADDR_WIDTH-1:61*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[62*CELL_ADDR_WIDTH-1:61*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[62*CELL_ADDR_WIDTH-1:61*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[62*CELL_ADDR_WIDTH-1:61*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[62*CELL_ADDR_WIDTH-1:61*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[62*CELL_ADDR_WIDTH-1:61*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_4_top[0])
				begin
				reg_FSM_to_Cell_read_addr[63*CELL_ADDR_WIDTH-1:62*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_top[1])
				begin
				reg_FSM_to_Cell_read_addr[63*CELL_ADDR_WIDTH-1:62*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_top[2])
				begin
				reg_FSM_to_Cell_read_addr[63*CELL_ADDR_WIDTH-1:62*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_top[3])
				begin
				reg_FSM_to_Cell_read_addr[63*CELL_ADDR_WIDTH-1:62*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_top[4])
				begin
				reg_FSM_to_Cell_read_addr[63*CELL_ADDR_WIDTH-1:62*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[63*CELL_ADDR_WIDTH-1:62*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[64*CELL_ADDR_WIDTH-1:63*CELL_ADDR_WIDTH] = 0;
			end
		3:
			begin
			reg_FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH] = 0;
			if (arbiter_1_1_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_1_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_1_top[0])
				begin
				reg_FSM_to_Cell_read_addr[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_top[1])
				begin
				reg_FSM_to_Cell_read_addr[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_top[2])
				begin
				reg_FSM_to_Cell_read_addr[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_top[3])
				begin
				reg_FSM_to_Cell_read_addr[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_top[4])
				begin
				reg_FSM_to_Cell_read_addr[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH] = 0;
			if (arbiter_1_2_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_2_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_2_top[0])
				begin
				reg_FSM_to_Cell_read_addr[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_top[1])
				begin
				reg_FSM_to_Cell_read_addr[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_top[2])
				begin
				reg_FSM_to_Cell_read_addr[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_top[3])
				begin
				reg_FSM_to_Cell_read_addr[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_top[4])
				begin
				reg_FSM_to_Cell_read_addr[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH] = 0;
			if (arbiter_1_3_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_3_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_3_top[0])
				begin
				reg_FSM_to_Cell_read_addr[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_top[1])
				begin
				reg_FSM_to_Cell_read_addr[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_top[2])
				begin
				reg_FSM_to_Cell_read_addr[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_top[3])
				begin
				reg_FSM_to_Cell_read_addr[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_top[4])
				begin
				reg_FSM_to_Cell_read_addr[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH] = 0;
			if (arbiter_1_4_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_4_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[15*CELL_ADDR_WIDTH-1:14*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[15*CELL_ADDR_WIDTH-1:14*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[15*CELL_ADDR_WIDTH-1:14*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[15*CELL_ADDR_WIDTH-1:14*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[15*CELL_ADDR_WIDTH-1:14*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[15*CELL_ADDR_WIDTH-1:14*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_4_top[0])
				begin
				reg_FSM_to_Cell_read_addr[16*CELL_ADDR_WIDTH-1:15*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_top[1])
				begin
				reg_FSM_to_Cell_read_addr[16*CELL_ADDR_WIDTH-1:15*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_top[2])
				begin
				reg_FSM_to_Cell_read_addr[16*CELL_ADDR_WIDTH-1:15*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_top[3])
				begin
				reg_FSM_to_Cell_read_addr[16*CELL_ADDR_WIDTH-1:15*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_top[4])
				begin
				reg_FSM_to_Cell_read_addr[16*CELL_ADDR_WIDTH-1:15*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[16*CELL_ADDR_WIDTH-1:15*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[17*CELL_ADDR_WIDTH-1:16*CELL_ADDR_WIDTH] = 0;
			if (arbiter_2_1_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[18*CELL_ADDR_WIDTH-1:17*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[18*CELL_ADDR_WIDTH-1:17*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[18*CELL_ADDR_WIDTH-1:17*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[18*CELL_ADDR_WIDTH-1:17*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[18*CELL_ADDR_WIDTH-1:17*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_1_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[19*CELL_ADDR_WIDTH-1:18*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[19*CELL_ADDR_WIDTH-1:18*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[19*CELL_ADDR_WIDTH-1:18*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[19*CELL_ADDR_WIDTH-1:18*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[19*CELL_ADDR_WIDTH-1:18*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[19*CELL_ADDR_WIDTH-1:18*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_1_top[0])
				begin
				reg_FSM_to_Cell_read_addr[20*CELL_ADDR_WIDTH-1:19*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_top[1])
				begin
				reg_FSM_to_Cell_read_addr[20*CELL_ADDR_WIDTH-1:19*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_top[2])
				begin
				reg_FSM_to_Cell_read_addr[20*CELL_ADDR_WIDTH-1:19*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_top[3])
				begin
				reg_FSM_to_Cell_read_addr[20*CELL_ADDR_WIDTH-1:19*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_top[4])
				begin
				reg_FSM_to_Cell_read_addr[20*CELL_ADDR_WIDTH-1:19*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[20*CELL_ADDR_WIDTH-1:19*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[21*CELL_ADDR_WIDTH-1:20*CELL_ADDR_WIDTH] = 0;
			if (arbiter_2_2_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[22*CELL_ADDR_WIDTH-1:21*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[22*CELL_ADDR_WIDTH-1:21*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[22*CELL_ADDR_WIDTH-1:21*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[22*CELL_ADDR_WIDTH-1:21*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[22*CELL_ADDR_WIDTH-1:21*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_2_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[23*CELL_ADDR_WIDTH-1:22*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[23*CELL_ADDR_WIDTH-1:22*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[23*CELL_ADDR_WIDTH-1:22*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[23*CELL_ADDR_WIDTH-1:22*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[23*CELL_ADDR_WIDTH-1:22*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[23*CELL_ADDR_WIDTH-1:22*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_2_top[0])
				begin
				reg_FSM_to_Cell_read_addr[24*CELL_ADDR_WIDTH-1:23*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_top[1])
				begin
				reg_FSM_to_Cell_read_addr[24*CELL_ADDR_WIDTH-1:23*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_top[2])
				begin
				reg_FSM_to_Cell_read_addr[24*CELL_ADDR_WIDTH-1:23*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_top[3])
				begin
				reg_FSM_to_Cell_read_addr[24*CELL_ADDR_WIDTH-1:23*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_top[4])
				begin
				reg_FSM_to_Cell_read_addr[24*CELL_ADDR_WIDTH-1:23*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[24*CELL_ADDR_WIDTH-1:23*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[25*CELL_ADDR_WIDTH-1:24*CELL_ADDR_WIDTH] = 0;
			if (arbiter_2_3_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[26*CELL_ADDR_WIDTH-1:25*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[26*CELL_ADDR_WIDTH-1:25*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[26*CELL_ADDR_WIDTH-1:25*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[26*CELL_ADDR_WIDTH-1:25*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[26*CELL_ADDR_WIDTH-1:25*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_3_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[27*CELL_ADDR_WIDTH-1:26*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[27*CELL_ADDR_WIDTH-1:26*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[27*CELL_ADDR_WIDTH-1:26*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[27*CELL_ADDR_WIDTH-1:26*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[27*CELL_ADDR_WIDTH-1:26*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[27*CELL_ADDR_WIDTH-1:26*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_3_top[0])
				begin
				reg_FSM_to_Cell_read_addr[28*CELL_ADDR_WIDTH-1:27*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_top[1])
				begin
				reg_FSM_to_Cell_read_addr[28*CELL_ADDR_WIDTH-1:27*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_top[2])
				begin
				reg_FSM_to_Cell_read_addr[28*CELL_ADDR_WIDTH-1:27*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_top[3])
				begin
				reg_FSM_to_Cell_read_addr[28*CELL_ADDR_WIDTH-1:27*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_top[4])
				begin
				reg_FSM_to_Cell_read_addr[28*CELL_ADDR_WIDTH-1:27*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[28*CELL_ADDR_WIDTH-1:27*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[29*CELL_ADDR_WIDTH-1:28*CELL_ADDR_WIDTH] = 0;
			if (arbiter_2_4_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[30*CELL_ADDR_WIDTH-1:29*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[30*CELL_ADDR_WIDTH-1:29*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[30*CELL_ADDR_WIDTH-1:29*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[30*CELL_ADDR_WIDTH-1:29*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[30*CELL_ADDR_WIDTH-1:29*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_4_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[31*CELL_ADDR_WIDTH-1:30*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[31*CELL_ADDR_WIDTH-1:30*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[31*CELL_ADDR_WIDTH-1:30*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[31*CELL_ADDR_WIDTH-1:30*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[31*CELL_ADDR_WIDTH-1:30*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[31*CELL_ADDR_WIDTH-1:30*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_4_top[0])
				begin
				reg_FSM_to_Cell_read_addr[32*CELL_ADDR_WIDTH-1:31*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_top[1])
				begin
				reg_FSM_to_Cell_read_addr[32*CELL_ADDR_WIDTH-1:31*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_top[2])
				begin
				reg_FSM_to_Cell_read_addr[32*CELL_ADDR_WIDTH-1:31*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_top[3])
				begin
				reg_FSM_to_Cell_read_addr[32*CELL_ADDR_WIDTH-1:31*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_top[4])
				begin
				reg_FSM_to_Cell_read_addr[32*CELL_ADDR_WIDTH-1:31*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[32*CELL_ADDR_WIDTH-1:31*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[33*CELL_ADDR_WIDTH-1:32*CELL_ADDR_WIDTH] = 0;
			if (arbiter_3_1_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[34*CELL_ADDR_WIDTH-1:33*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[34*CELL_ADDR_WIDTH-1:33*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[34*CELL_ADDR_WIDTH-1:33*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[34*CELL_ADDR_WIDTH-1:33*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[34*CELL_ADDR_WIDTH-1:33*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_1_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[35*CELL_ADDR_WIDTH-1:34*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[35*CELL_ADDR_WIDTH-1:34*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[35*CELL_ADDR_WIDTH-1:34*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[35*CELL_ADDR_WIDTH-1:34*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[35*CELL_ADDR_WIDTH-1:34*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[35*CELL_ADDR_WIDTH-1:34*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_1_top[0])
				begin
				reg_FSM_to_Cell_read_addr[36*CELL_ADDR_WIDTH-1:35*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_top[1])
				begin
				reg_FSM_to_Cell_read_addr[36*CELL_ADDR_WIDTH-1:35*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_top[2])
				begin
				reg_FSM_to_Cell_read_addr[36*CELL_ADDR_WIDTH-1:35*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_top[3])
				begin
				reg_FSM_to_Cell_read_addr[36*CELL_ADDR_WIDTH-1:35*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_top[4])
				begin
				reg_FSM_to_Cell_read_addr[36*CELL_ADDR_WIDTH-1:35*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[36*CELL_ADDR_WIDTH-1:35*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[37*CELL_ADDR_WIDTH-1:36*CELL_ADDR_WIDTH] = 0;
			if (arbiter_3_2_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[38*CELL_ADDR_WIDTH-1:37*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[38*CELL_ADDR_WIDTH-1:37*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[38*CELL_ADDR_WIDTH-1:37*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[38*CELL_ADDR_WIDTH-1:37*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[38*CELL_ADDR_WIDTH-1:37*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_2_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[39*CELL_ADDR_WIDTH-1:38*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[39*CELL_ADDR_WIDTH-1:38*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[39*CELL_ADDR_WIDTH-1:38*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[39*CELL_ADDR_WIDTH-1:38*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[39*CELL_ADDR_WIDTH-1:38*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[39*CELL_ADDR_WIDTH-1:38*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_2_top[0])
				begin
				reg_FSM_to_Cell_read_addr[40*CELL_ADDR_WIDTH-1:39*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_top[1])
				begin
				reg_FSM_to_Cell_read_addr[40*CELL_ADDR_WIDTH-1:39*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_top[2])
				begin
				reg_FSM_to_Cell_read_addr[40*CELL_ADDR_WIDTH-1:39*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_top[3])
				begin
				reg_FSM_to_Cell_read_addr[40*CELL_ADDR_WIDTH-1:39*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_top[4])
				begin
				reg_FSM_to_Cell_read_addr[40*CELL_ADDR_WIDTH-1:39*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[40*CELL_ADDR_WIDTH-1:39*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[41*CELL_ADDR_WIDTH-1:40*CELL_ADDR_WIDTH] = 0;
			if (arbiter_3_3_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[42*CELL_ADDR_WIDTH-1:41*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[42*CELL_ADDR_WIDTH-1:41*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[42*CELL_ADDR_WIDTH-1:41*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[42*CELL_ADDR_WIDTH-1:41*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[42*CELL_ADDR_WIDTH-1:41*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_3_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[43*CELL_ADDR_WIDTH-1:42*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[43*CELL_ADDR_WIDTH-1:42*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[43*CELL_ADDR_WIDTH-1:42*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[43*CELL_ADDR_WIDTH-1:42*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[43*CELL_ADDR_WIDTH-1:42*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[43*CELL_ADDR_WIDTH-1:42*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_3_top[0])
				begin
				reg_FSM_to_Cell_read_addr[44*CELL_ADDR_WIDTH-1:43*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_top[1])
				begin
				reg_FSM_to_Cell_read_addr[44*CELL_ADDR_WIDTH-1:43*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_top[2])
				begin
				reg_FSM_to_Cell_read_addr[44*CELL_ADDR_WIDTH-1:43*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_top[3])
				begin
				reg_FSM_to_Cell_read_addr[44*CELL_ADDR_WIDTH-1:43*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_top[4])
				begin
				reg_FSM_to_Cell_read_addr[44*CELL_ADDR_WIDTH-1:43*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[44*CELL_ADDR_WIDTH-1:43*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[45*CELL_ADDR_WIDTH-1:44*CELL_ADDR_WIDTH] = 0;
			if (arbiter_3_4_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[46*CELL_ADDR_WIDTH-1:45*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[46*CELL_ADDR_WIDTH-1:45*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[46*CELL_ADDR_WIDTH-1:45*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[46*CELL_ADDR_WIDTH-1:45*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[46*CELL_ADDR_WIDTH-1:45*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_4_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[47*CELL_ADDR_WIDTH-1:46*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[47*CELL_ADDR_WIDTH-1:46*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[47*CELL_ADDR_WIDTH-1:46*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[47*CELL_ADDR_WIDTH-1:46*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[47*CELL_ADDR_WIDTH-1:46*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[47*CELL_ADDR_WIDTH-1:46*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_4_top[0])
				begin
				reg_FSM_to_Cell_read_addr[48*CELL_ADDR_WIDTH-1:47*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_top[1])
				begin
				reg_FSM_to_Cell_read_addr[48*CELL_ADDR_WIDTH-1:47*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_top[2])
				begin
				reg_FSM_to_Cell_read_addr[48*CELL_ADDR_WIDTH-1:47*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_top[3])
				begin
				reg_FSM_to_Cell_read_addr[48*CELL_ADDR_WIDTH-1:47*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_top[4])
				begin
				reg_FSM_to_Cell_read_addr[48*CELL_ADDR_WIDTH-1:47*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[48*CELL_ADDR_WIDTH-1:47*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[49*CELL_ADDR_WIDTH-1:48*CELL_ADDR_WIDTH] = 0;
			if (arbiter_4_1_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[50*CELL_ADDR_WIDTH-1:49*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[50*CELL_ADDR_WIDTH-1:49*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[50*CELL_ADDR_WIDTH-1:49*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[50*CELL_ADDR_WIDTH-1:49*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[50*CELL_ADDR_WIDTH-1:49*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_1_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[51*CELL_ADDR_WIDTH-1:50*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[51*CELL_ADDR_WIDTH-1:50*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[51*CELL_ADDR_WIDTH-1:50*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[51*CELL_ADDR_WIDTH-1:50*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[51*CELL_ADDR_WIDTH-1:50*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[51*CELL_ADDR_WIDTH-1:50*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_1_top[0])
				begin
				reg_FSM_to_Cell_read_addr[52*CELL_ADDR_WIDTH-1:51*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_top[1])
				begin
				reg_FSM_to_Cell_read_addr[52*CELL_ADDR_WIDTH-1:51*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_top[2])
				begin
				reg_FSM_to_Cell_read_addr[52*CELL_ADDR_WIDTH-1:51*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_top[3])
				begin
				reg_FSM_to_Cell_read_addr[52*CELL_ADDR_WIDTH-1:51*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_top[4])
				begin
				reg_FSM_to_Cell_read_addr[52*CELL_ADDR_WIDTH-1:51*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[52*CELL_ADDR_WIDTH-1:51*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[53*CELL_ADDR_WIDTH-1:52*CELL_ADDR_WIDTH] = 0;
			if (arbiter_4_2_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[54*CELL_ADDR_WIDTH-1:53*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[54*CELL_ADDR_WIDTH-1:53*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[54*CELL_ADDR_WIDTH-1:53*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[54*CELL_ADDR_WIDTH-1:53*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[54*CELL_ADDR_WIDTH-1:53*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_2_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[55*CELL_ADDR_WIDTH-1:54*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[55*CELL_ADDR_WIDTH-1:54*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[55*CELL_ADDR_WIDTH-1:54*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[55*CELL_ADDR_WIDTH-1:54*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[55*CELL_ADDR_WIDTH-1:54*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[55*CELL_ADDR_WIDTH-1:54*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_2_top[0])
				begin
				reg_FSM_to_Cell_read_addr[56*CELL_ADDR_WIDTH-1:55*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_top[1])
				begin
				reg_FSM_to_Cell_read_addr[56*CELL_ADDR_WIDTH-1:55*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_top[2])
				begin
				reg_FSM_to_Cell_read_addr[56*CELL_ADDR_WIDTH-1:55*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_top[3])
				begin
				reg_FSM_to_Cell_read_addr[56*CELL_ADDR_WIDTH-1:55*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_top[4])
				begin
				reg_FSM_to_Cell_read_addr[56*CELL_ADDR_WIDTH-1:55*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[56*CELL_ADDR_WIDTH-1:55*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[57*CELL_ADDR_WIDTH-1:56*CELL_ADDR_WIDTH] = 0;
			if (arbiter_4_3_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[58*CELL_ADDR_WIDTH-1:57*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[58*CELL_ADDR_WIDTH-1:57*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[58*CELL_ADDR_WIDTH-1:57*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[58*CELL_ADDR_WIDTH-1:57*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[58*CELL_ADDR_WIDTH-1:57*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_3_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[59*CELL_ADDR_WIDTH-1:58*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[59*CELL_ADDR_WIDTH-1:58*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[59*CELL_ADDR_WIDTH-1:58*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[59*CELL_ADDR_WIDTH-1:58*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[59*CELL_ADDR_WIDTH-1:58*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[59*CELL_ADDR_WIDTH-1:58*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_3_top[0])
				begin
				reg_FSM_to_Cell_read_addr[60*CELL_ADDR_WIDTH-1:59*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_top[1])
				begin
				reg_FSM_to_Cell_read_addr[60*CELL_ADDR_WIDTH-1:59*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_top[2])
				begin
				reg_FSM_to_Cell_read_addr[60*CELL_ADDR_WIDTH-1:59*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_top[3])
				begin
				reg_FSM_to_Cell_read_addr[60*CELL_ADDR_WIDTH-1:59*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_top[4])
				begin
				reg_FSM_to_Cell_read_addr[60*CELL_ADDR_WIDTH-1:59*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[60*CELL_ADDR_WIDTH-1:59*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[61*CELL_ADDR_WIDTH-1:60*CELL_ADDR_WIDTH] = 0;
			if (arbiter_4_4_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[62*CELL_ADDR_WIDTH-1:61*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[62*CELL_ADDR_WIDTH-1:61*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[62*CELL_ADDR_WIDTH-1:61*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[62*CELL_ADDR_WIDTH-1:61*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[62*CELL_ADDR_WIDTH-1:61*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_4_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[63*CELL_ADDR_WIDTH-1:62*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[63*CELL_ADDR_WIDTH-1:62*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[63*CELL_ADDR_WIDTH-1:62*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[63*CELL_ADDR_WIDTH-1:62*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[63*CELL_ADDR_WIDTH-1:62*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[63*CELL_ADDR_WIDTH-1:62*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_4_top[0])
				begin
				reg_FSM_to_Cell_read_addr[64*CELL_ADDR_WIDTH-1:63*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_top[1])
				begin
				reg_FSM_to_Cell_read_addr[64*CELL_ADDR_WIDTH-1:63*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_top[2])
				begin
				reg_FSM_to_Cell_read_addr[64*CELL_ADDR_WIDTH-1:63*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_top[3])
				begin
				reg_FSM_to_Cell_read_addr[64*CELL_ADDR_WIDTH-1:63*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_top[4])
				begin
				reg_FSM_to_Cell_read_addr[64*CELL_ADDR_WIDTH-1:63*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[64*CELL_ADDR_WIDTH-1:63*CELL_ADDR_WIDTH] = 0;
				end
			end
		4:
			begin
			if (arbiter_1_1_top[0])
				begin
				reg_FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_top[1])
				begin
				reg_FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_top[2])
				begin
				reg_FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_top[3])
				begin
				reg_FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_top[4])
				begin
				reg_FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH] = 0;
			if (arbiter_1_1_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_1_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_1_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_2_top[0])
				begin
				reg_FSM_to_Cell_read_addr[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_top[1])
				begin
				reg_FSM_to_Cell_read_addr[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_top[2])
				begin
				reg_FSM_to_Cell_read_addr[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_top[3])
				begin
				reg_FSM_to_Cell_read_addr[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_top[4])
				begin
				reg_FSM_to_Cell_read_addr[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH] = 0;
			if (arbiter_1_2_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_2_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_2_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_3_top[0])
				begin
				reg_FSM_to_Cell_read_addr[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_top[1])
				begin
				reg_FSM_to_Cell_read_addr[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_top[2])
				begin
				reg_FSM_to_Cell_read_addr[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_top[3])
				begin
				reg_FSM_to_Cell_read_addr[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_top[4])
				begin
				reg_FSM_to_Cell_read_addr[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH] = 0;
			if (arbiter_1_3_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_3_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_3_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_4_top[0])
				begin
				reg_FSM_to_Cell_read_addr[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_top[1])
				begin
				reg_FSM_to_Cell_read_addr[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_top[2])
				begin
				reg_FSM_to_Cell_read_addr[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_top[3])
				begin
				reg_FSM_to_Cell_read_addr[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_top[4])
				begin
				reg_FSM_to_Cell_read_addr[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH] = 0;
			if (arbiter_1_4_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[15*CELL_ADDR_WIDTH-1:14*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[15*CELL_ADDR_WIDTH-1:14*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[15*CELL_ADDR_WIDTH-1:14*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[15*CELL_ADDR_WIDTH-1:14*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[15*CELL_ADDR_WIDTH-1:14*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_1_4_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[16*CELL_ADDR_WIDTH-1:15*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[16*CELL_ADDR_WIDTH-1:15*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[16*CELL_ADDR_WIDTH-1:15*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[16*CELL_ADDR_WIDTH-1:15*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_1_4_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[16*CELL_ADDR_WIDTH-1:15*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[16*CELL_ADDR_WIDTH-1:15*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_1_top[0])
				begin
				reg_FSM_to_Cell_read_addr[17*CELL_ADDR_WIDTH-1:16*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_top[1])
				begin
				reg_FSM_to_Cell_read_addr[17*CELL_ADDR_WIDTH-1:16*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_top[2])
				begin
				reg_FSM_to_Cell_read_addr[17*CELL_ADDR_WIDTH-1:16*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_top[3])
				begin
				reg_FSM_to_Cell_read_addr[17*CELL_ADDR_WIDTH-1:16*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_top[4])
				begin
				reg_FSM_to_Cell_read_addr[17*CELL_ADDR_WIDTH-1:16*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[17*CELL_ADDR_WIDTH-1:16*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[18*CELL_ADDR_WIDTH-1:17*CELL_ADDR_WIDTH] = 0;
			if (arbiter_2_1_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[19*CELL_ADDR_WIDTH-1:18*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[19*CELL_ADDR_WIDTH-1:18*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[19*CELL_ADDR_WIDTH-1:18*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[19*CELL_ADDR_WIDTH-1:18*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[19*CELL_ADDR_WIDTH-1:18*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_1_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[20*CELL_ADDR_WIDTH-1:19*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[20*CELL_ADDR_WIDTH-1:19*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[20*CELL_ADDR_WIDTH-1:19*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[20*CELL_ADDR_WIDTH-1:19*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_1_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[20*CELL_ADDR_WIDTH-1:19*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[20*CELL_ADDR_WIDTH-1:19*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_2_top[0])
				begin
				reg_FSM_to_Cell_read_addr[21*CELL_ADDR_WIDTH-1:20*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_top[1])
				begin
				reg_FSM_to_Cell_read_addr[21*CELL_ADDR_WIDTH-1:20*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_top[2])
				begin
				reg_FSM_to_Cell_read_addr[21*CELL_ADDR_WIDTH-1:20*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_top[3])
				begin
				reg_FSM_to_Cell_read_addr[21*CELL_ADDR_WIDTH-1:20*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_top[4])
				begin
				reg_FSM_to_Cell_read_addr[21*CELL_ADDR_WIDTH-1:20*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[21*CELL_ADDR_WIDTH-1:20*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[22*CELL_ADDR_WIDTH-1:21*CELL_ADDR_WIDTH] = 0;
			if (arbiter_2_2_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[23*CELL_ADDR_WIDTH-1:22*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[23*CELL_ADDR_WIDTH-1:22*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[23*CELL_ADDR_WIDTH-1:22*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[23*CELL_ADDR_WIDTH-1:22*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[23*CELL_ADDR_WIDTH-1:22*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_2_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[24*CELL_ADDR_WIDTH-1:23*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[24*CELL_ADDR_WIDTH-1:23*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[24*CELL_ADDR_WIDTH-1:23*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[24*CELL_ADDR_WIDTH-1:23*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_2_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[24*CELL_ADDR_WIDTH-1:23*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[24*CELL_ADDR_WIDTH-1:23*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_3_top[0])
				begin
				reg_FSM_to_Cell_read_addr[25*CELL_ADDR_WIDTH-1:24*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_top[1])
				begin
				reg_FSM_to_Cell_read_addr[25*CELL_ADDR_WIDTH-1:24*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_top[2])
				begin
				reg_FSM_to_Cell_read_addr[25*CELL_ADDR_WIDTH-1:24*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_top[3])
				begin
				reg_FSM_to_Cell_read_addr[25*CELL_ADDR_WIDTH-1:24*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_top[4])
				begin
				reg_FSM_to_Cell_read_addr[25*CELL_ADDR_WIDTH-1:24*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[25*CELL_ADDR_WIDTH-1:24*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[26*CELL_ADDR_WIDTH-1:25*CELL_ADDR_WIDTH] = 0;
			if (arbiter_2_3_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[27*CELL_ADDR_WIDTH-1:26*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[27*CELL_ADDR_WIDTH-1:26*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[27*CELL_ADDR_WIDTH-1:26*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[27*CELL_ADDR_WIDTH-1:26*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[27*CELL_ADDR_WIDTH-1:26*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_3_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[28*CELL_ADDR_WIDTH-1:27*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_2[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[28*CELL_ADDR_WIDTH-1:27*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[28*CELL_ADDR_WIDTH-1:27*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[28*CELL_ADDR_WIDTH-1:27*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_3_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[28*CELL_ADDR_WIDTH-1:27*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[28*CELL_ADDR_WIDTH-1:27*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_4_top[0])
				begin
				reg_FSM_to_Cell_read_addr[29*CELL_ADDR_WIDTH-1:28*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_top[1])
				begin
				reg_FSM_to_Cell_read_addr[29*CELL_ADDR_WIDTH-1:28*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_top[2])
				begin
				reg_FSM_to_Cell_read_addr[29*CELL_ADDR_WIDTH-1:28*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_top[3])
				begin
				reg_FSM_to_Cell_read_addr[29*CELL_ADDR_WIDTH-1:28*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_top[4])
				begin
				reg_FSM_to_Cell_read_addr[29*CELL_ADDR_WIDTH-1:28*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[29*CELL_ADDR_WIDTH-1:28*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[30*CELL_ADDR_WIDTH-1:29*CELL_ADDR_WIDTH] = 0;
			if (arbiter_2_4_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[31*CELL_ADDR_WIDTH-1:30*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[31*CELL_ADDR_WIDTH-1:30*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[31*CELL_ADDR_WIDTH-1:30*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[31*CELL_ADDR_WIDTH-1:30*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[31*CELL_ADDR_WIDTH-1:30*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_2_4_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[32*CELL_ADDR_WIDTH-1:31*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_1[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[32*CELL_ADDR_WIDTH-1:31*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_3[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[32*CELL_ADDR_WIDTH-1:31*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_1_4[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[32*CELL_ADDR_WIDTH-1:31*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_2_4_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[32*CELL_ADDR_WIDTH-1:31*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[32*CELL_ADDR_WIDTH-1:31*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_1_top[0])
				begin
				reg_FSM_to_Cell_read_addr[33*CELL_ADDR_WIDTH-1:32*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_top[1])
				begin
				reg_FSM_to_Cell_read_addr[33*CELL_ADDR_WIDTH-1:32*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_top[2])
				begin
				reg_FSM_to_Cell_read_addr[33*CELL_ADDR_WIDTH-1:32*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_top[3])
				begin
				reg_FSM_to_Cell_read_addr[33*CELL_ADDR_WIDTH-1:32*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_top[4])
				begin
				reg_FSM_to_Cell_read_addr[33*CELL_ADDR_WIDTH-1:32*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[33*CELL_ADDR_WIDTH-1:32*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[34*CELL_ADDR_WIDTH-1:33*CELL_ADDR_WIDTH] = 0;
			if (arbiter_3_1_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[35*CELL_ADDR_WIDTH-1:34*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[35*CELL_ADDR_WIDTH-1:34*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[35*CELL_ADDR_WIDTH-1:34*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[35*CELL_ADDR_WIDTH-1:34*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[35*CELL_ADDR_WIDTH-1:34*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_1_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[36*CELL_ADDR_WIDTH-1:35*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[36*CELL_ADDR_WIDTH-1:35*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[36*CELL_ADDR_WIDTH-1:35*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[36*CELL_ADDR_WIDTH-1:35*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_1_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[36*CELL_ADDR_WIDTH-1:35*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[36*CELL_ADDR_WIDTH-1:35*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_2_top[0])
				begin
				reg_FSM_to_Cell_read_addr[37*CELL_ADDR_WIDTH-1:36*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_top[1])
				begin
				reg_FSM_to_Cell_read_addr[37*CELL_ADDR_WIDTH-1:36*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_top[2])
				begin
				reg_FSM_to_Cell_read_addr[37*CELL_ADDR_WIDTH-1:36*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_top[3])
				begin
				reg_FSM_to_Cell_read_addr[37*CELL_ADDR_WIDTH-1:36*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_top[4])
				begin
				reg_FSM_to_Cell_read_addr[37*CELL_ADDR_WIDTH-1:36*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[37*CELL_ADDR_WIDTH-1:36*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[38*CELL_ADDR_WIDTH-1:37*CELL_ADDR_WIDTH] = 0;
			if (arbiter_3_2_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[39*CELL_ADDR_WIDTH-1:38*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[39*CELL_ADDR_WIDTH-1:38*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[39*CELL_ADDR_WIDTH-1:38*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[39*CELL_ADDR_WIDTH-1:38*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[39*CELL_ADDR_WIDTH-1:38*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_2_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[40*CELL_ADDR_WIDTH-1:39*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[40*CELL_ADDR_WIDTH-1:39*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[40*CELL_ADDR_WIDTH-1:39*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[40*CELL_ADDR_WIDTH-1:39*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_2_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[40*CELL_ADDR_WIDTH-1:39*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[40*CELL_ADDR_WIDTH-1:39*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_3_top[0])
				begin
				reg_FSM_to_Cell_read_addr[41*CELL_ADDR_WIDTH-1:40*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_top[1])
				begin
				reg_FSM_to_Cell_read_addr[41*CELL_ADDR_WIDTH-1:40*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_top[2])
				begin
				reg_FSM_to_Cell_read_addr[41*CELL_ADDR_WIDTH-1:40*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_top[3])
				begin
				reg_FSM_to_Cell_read_addr[41*CELL_ADDR_WIDTH-1:40*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_top[4])
				begin
				reg_FSM_to_Cell_read_addr[41*CELL_ADDR_WIDTH-1:40*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[41*CELL_ADDR_WIDTH-1:40*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[42*CELL_ADDR_WIDTH-1:41*CELL_ADDR_WIDTH] = 0;
			if (arbiter_3_3_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[43*CELL_ADDR_WIDTH-1:42*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[43*CELL_ADDR_WIDTH-1:42*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[43*CELL_ADDR_WIDTH-1:42*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[43*CELL_ADDR_WIDTH-1:42*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[43*CELL_ADDR_WIDTH-1:42*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_3_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[44*CELL_ADDR_WIDTH-1:43*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_2[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[44*CELL_ADDR_WIDTH-1:43*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[44*CELL_ADDR_WIDTH-1:43*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[44*CELL_ADDR_WIDTH-1:43*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_3_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[44*CELL_ADDR_WIDTH-1:43*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[44*CELL_ADDR_WIDTH-1:43*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_4_top[0])
				begin
				reg_FSM_to_Cell_read_addr[45*CELL_ADDR_WIDTH-1:44*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_top[1])
				begin
				reg_FSM_to_Cell_read_addr[45*CELL_ADDR_WIDTH-1:44*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_top[2])
				begin
				reg_FSM_to_Cell_read_addr[45*CELL_ADDR_WIDTH-1:44*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_top[3])
				begin
				reg_FSM_to_Cell_read_addr[45*CELL_ADDR_WIDTH-1:44*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_top[4])
				begin
				reg_FSM_to_Cell_read_addr[45*CELL_ADDR_WIDTH-1:44*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[45*CELL_ADDR_WIDTH-1:44*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[46*CELL_ADDR_WIDTH-1:45*CELL_ADDR_WIDTH] = 0;
			if (arbiter_3_4_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[47*CELL_ADDR_WIDTH-1:46*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[47*CELL_ADDR_WIDTH-1:46*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[47*CELL_ADDR_WIDTH-1:46*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[47*CELL_ADDR_WIDTH-1:46*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[47*CELL_ADDR_WIDTH-1:46*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_3_4_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[48*CELL_ADDR_WIDTH-1:47*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_1[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[48*CELL_ADDR_WIDTH-1:47*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_3[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[48*CELL_ADDR_WIDTH-1:47*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_2_4[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[48*CELL_ADDR_WIDTH-1:47*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_3_4_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[48*CELL_ADDR_WIDTH-1:47*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[48*CELL_ADDR_WIDTH-1:47*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_1_top[0])
				begin
				reg_FSM_to_Cell_read_addr[49*CELL_ADDR_WIDTH-1:48*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_top[1])
				begin
				reg_FSM_to_Cell_read_addr[49*CELL_ADDR_WIDTH-1:48*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_top[2])
				begin
				reg_FSM_to_Cell_read_addr[49*CELL_ADDR_WIDTH-1:48*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_top[3])
				begin
				reg_FSM_to_Cell_read_addr[49*CELL_ADDR_WIDTH-1:48*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_top[4])
				begin
				reg_FSM_to_Cell_read_addr[49*CELL_ADDR_WIDTH-1:48*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[49*CELL_ADDR_WIDTH-1:48*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[50*CELL_ADDR_WIDTH-1:49*CELL_ADDR_WIDTH] = 0;
			if (arbiter_4_1_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[51*CELL_ADDR_WIDTH-1:50*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[51*CELL_ADDR_WIDTH-1:50*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[51*CELL_ADDR_WIDTH-1:50*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[51*CELL_ADDR_WIDTH-1:50*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[51*CELL_ADDR_WIDTH-1:50*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_1_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[52*CELL_ADDR_WIDTH-1:51*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[52*CELL_ADDR_WIDTH-1:51*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[52*CELL_ADDR_WIDTH-1:51*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[52*CELL_ADDR_WIDTH-1:51*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_1_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[52*CELL_ADDR_WIDTH-1:51*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[52*CELL_ADDR_WIDTH-1:51*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_2_top[0])
				begin
				reg_FSM_to_Cell_read_addr[53*CELL_ADDR_WIDTH-1:52*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_top[1])
				begin
				reg_FSM_to_Cell_read_addr[53*CELL_ADDR_WIDTH-1:52*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_top[2])
				begin
				reg_FSM_to_Cell_read_addr[53*CELL_ADDR_WIDTH-1:52*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_top[3])
				begin
				reg_FSM_to_Cell_read_addr[53*CELL_ADDR_WIDTH-1:52*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_top[4])
				begin
				reg_FSM_to_Cell_read_addr[53*CELL_ADDR_WIDTH-1:52*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[53*CELL_ADDR_WIDTH-1:52*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[54*CELL_ADDR_WIDTH-1:53*CELL_ADDR_WIDTH] = 0;
			if (arbiter_4_2_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[55*CELL_ADDR_WIDTH-1:54*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[55*CELL_ADDR_WIDTH-1:54*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[55*CELL_ADDR_WIDTH-1:54*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[55*CELL_ADDR_WIDTH-1:54*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[55*CELL_ADDR_WIDTH-1:54*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_2_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[56*CELL_ADDR_WIDTH-1:55*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[56*CELL_ADDR_WIDTH-1:55*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[56*CELL_ADDR_WIDTH-1:55*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[56*CELL_ADDR_WIDTH-1:55*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_1[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_2_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[56*CELL_ADDR_WIDTH-1:55*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[56*CELL_ADDR_WIDTH-1:55*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_3_top[0])
				begin
				reg_FSM_to_Cell_read_addr[57*CELL_ADDR_WIDTH-1:56*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_top[1])
				begin
				reg_FSM_to_Cell_read_addr[57*CELL_ADDR_WIDTH-1:56*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_top[2])
				begin
				reg_FSM_to_Cell_read_addr[57*CELL_ADDR_WIDTH-1:56*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_top[3])
				begin
				reg_FSM_to_Cell_read_addr[57*CELL_ADDR_WIDTH-1:56*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_top[4])
				begin
				reg_FSM_to_Cell_read_addr[57*CELL_ADDR_WIDTH-1:56*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[57*CELL_ADDR_WIDTH-1:56*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[58*CELL_ADDR_WIDTH-1:57*CELL_ADDR_WIDTH] = 0;
			if (arbiter_4_3_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[59*CELL_ADDR_WIDTH-1:58*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[59*CELL_ADDR_WIDTH-1:58*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[59*CELL_ADDR_WIDTH-1:58*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[59*CELL_ADDR_WIDTH-1:58*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[59*CELL_ADDR_WIDTH-1:58*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_3_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[60*CELL_ADDR_WIDTH-1:59*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_2[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[60*CELL_ADDR_WIDTH-1:59*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[60*CELL_ADDR_WIDTH-1:59*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[60*CELL_ADDR_WIDTH-1:59*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_2[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_3_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[60*CELL_ADDR_WIDTH-1:59*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[60*CELL_ADDR_WIDTH-1:59*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_4_top[0])
				begin
				reg_FSM_to_Cell_read_addr[61*CELL_ADDR_WIDTH-1:60*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_top[1])
				begin
				reg_FSM_to_Cell_read_addr[61*CELL_ADDR_WIDTH-1:60*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_top[2])
				begin
				reg_FSM_to_Cell_read_addr[61*CELL_ADDR_WIDTH-1:60*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_top[3])
				begin
				reg_FSM_to_Cell_read_addr[61*CELL_ADDR_WIDTH-1:60*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_top[4])
				begin
				reg_FSM_to_Cell_read_addr[61*CELL_ADDR_WIDTH-1:60*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[61*CELL_ADDR_WIDTH-1:60*CELL_ADDR_WIDTH] = 0;
				end
			reg_FSM_to_Cell_read_addr[62*CELL_ADDR_WIDTH-1:61*CELL_ADDR_WIDTH] = 0;
			if (arbiter_4_4_bottom[0])
				begin
				reg_FSM_to_Cell_read_addr[63*CELL_ADDR_WIDTH-1:62*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_bottom[1])
				begin
				reg_FSM_to_Cell_read_addr[63*CELL_ADDR_WIDTH-1:62*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_bottom[2])
				begin
				reg_FSM_to_Cell_read_addr[63*CELL_ADDR_WIDTH-1:62*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_bottom[3])
				begin
				reg_FSM_to_Cell_read_addr[63*CELL_ADDR_WIDTH-1:62*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[63*CELL_ADDR_WIDTH-1:62*CELL_ADDR_WIDTH] = 0;
				end
			if (arbiter_4_4_mid[0])
				begin
				reg_FSM_to_Cell_read_addr[64*CELL_ADDR_WIDTH-1:63*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_1[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_mid[1])
				begin
				reg_FSM_to_Cell_read_addr[64*CELL_ADDR_WIDTH-1:63*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_3[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_mid[2])
				begin
				reg_FSM_to_Cell_read_addr[64*CELL_ADDR_WIDTH-1:63*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_3_4[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_mid[3])
				begin
				reg_FSM_to_Cell_read_addr[64*CELL_ADDR_WIDTH-1:63*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_3[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				end
			else if (arbiter_4_4_mid[4])
				begin
				reg_FSM_to_Cell_read_addr[64*CELL_ADDR_WIDTH-1:63*CELL_ADDR_WIDTH] = FSM_to_Cell_read_addr_4_4[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				end
			else
				begin
				reg_FSM_to_Cell_read_addr[64*CELL_ADDR_WIDTH-1:63*CELL_ADDR_WIDTH] = 0;
				end
			end
		default:
			begin
			reg_FSM_to_Cell_read_addr = 0;
			end
	endcase
	reg_Cell_to_FSM_read_success_bit_1_1[0] = (arbiter_1_1_mid[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_4[3] = (arbiter_1_1_mid[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_1[9] = (arbiter_1_1_mid[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_2[6] = (arbiter_1_1_mid[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_4[12] = (arbiter_1_1_mid[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_1[1] = (arbiter_1_1_top[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_4[4] = (arbiter_1_1_top[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_1[10] = (arbiter_1_1_top[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_2[7] = (arbiter_1_1_top[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_4[13] = (arbiter_1_1_top[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_4[2] = (arbiter_1_1_bottom[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_1[8] = (arbiter_1_1_bottom[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_2[5] = (arbiter_1_1_bottom[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_4[11] = (arbiter_1_1_bottom[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_1[3] = (arbiter_1_2_mid[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_2[0] = (arbiter_1_2_mid[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_1[12] = (arbiter_1_2_mid[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_2[9] = (arbiter_1_2_mid[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_3[6] = (arbiter_1_2_mid[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_1[4] = (arbiter_1_2_top[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_2[1] = (arbiter_1_2_top[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_1[13] = (arbiter_1_2_top[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_2[10] = (arbiter_1_2_top[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_3[7] = (arbiter_1_2_top[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_1[2] = (arbiter_1_2_bottom[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_1[11] = (arbiter_1_2_bottom[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_2[8] = (arbiter_1_2_bottom[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_3[5] = (arbiter_1_2_bottom[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_2[3] = (arbiter_1_3_mid[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_3[0] = (arbiter_1_3_mid[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_2[12] = (arbiter_1_3_mid[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_3[9] = (arbiter_1_3_mid[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_4[6] = (arbiter_1_3_mid[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_2[4] = (arbiter_1_3_top[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_3[1] = (arbiter_1_3_top[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_2[13] = (arbiter_1_3_top[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_3[10] = (arbiter_1_3_top[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_4[7] = (arbiter_1_3_top[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_2[2] = (arbiter_1_3_bottom[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_2[11] = (arbiter_1_3_bottom[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_3[8] = (arbiter_1_3_bottom[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_4[5] = (arbiter_1_3_bottom[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_3[3] = (arbiter_1_4_mid[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_4[0] = (arbiter_1_4_mid[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_1[6] = (arbiter_1_4_mid[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_3[12] = (arbiter_1_4_mid[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_4[9] = (arbiter_1_4_mid[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_3[4] = (arbiter_1_4_top[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_4[1] = (arbiter_1_4_top[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_1[7] = (arbiter_1_4_top[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_3[13] = (arbiter_1_4_top[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_4[10] = (arbiter_1_4_top[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_3[2] = (arbiter_1_4_bottom[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_1[5] = (arbiter_1_4_bottom[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_3[11] = (arbiter_1_4_bottom[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_4[8] = (arbiter_1_4_bottom[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_1[9] = (arbiter_2_1_mid[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_2[6] = (arbiter_2_1_mid[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_4[12] = (arbiter_2_1_mid[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_1[0] = (arbiter_2_1_mid[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_4[3] = (arbiter_2_1_mid[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_1[10] = (arbiter_2_1_top[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_2[7] = (arbiter_2_1_top[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_4[13] = (arbiter_2_1_top[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_1[1] = (arbiter_2_1_top[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_4[4] = (arbiter_2_1_top[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_1[8] = (arbiter_2_1_bottom[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_2[5] = (arbiter_2_1_bottom[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_4[11] = (arbiter_2_1_bottom[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_4[2] = (arbiter_2_1_bottom[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_1[12] = (arbiter_2_2_mid[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_2[9] = (arbiter_2_2_mid[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_3[6] = (arbiter_2_2_mid[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_1[3] = (arbiter_2_2_mid[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_2[0] = (arbiter_2_2_mid[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_1[13] = (arbiter_2_2_top[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_2[10] = (arbiter_2_2_top[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_3[7] = (arbiter_2_2_top[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_1[4] = (arbiter_2_2_top[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_2[1] = (arbiter_2_2_top[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_1[11] = (arbiter_2_2_bottom[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_2[8] = (arbiter_2_2_bottom[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_3[5] = (arbiter_2_2_bottom[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_1[2] = (arbiter_2_2_bottom[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_2[12] = (arbiter_2_3_mid[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_3[9] = (arbiter_2_3_mid[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_4[6] = (arbiter_2_3_mid[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_2[3] = (arbiter_2_3_mid[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_3[0] = (arbiter_2_3_mid[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_2[13] = (arbiter_2_3_top[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_3[10] = (arbiter_2_3_top[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_4[7] = (arbiter_2_3_top[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_2[4] = (arbiter_2_3_top[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_3[1] = (arbiter_2_3_top[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_2[11] = (arbiter_2_3_bottom[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_3[8] = (arbiter_2_3_bottom[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_4[5] = (arbiter_2_3_bottom[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_2[2] = (arbiter_2_3_bottom[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_1[6] = (arbiter_2_4_mid[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_3[12] = (arbiter_2_4_mid[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_4[9] = (arbiter_2_4_mid[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_3[3] = (arbiter_2_4_mid[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_4[0] = (arbiter_2_4_mid[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_1[7] = (arbiter_2_4_top[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_3[13] = (arbiter_2_4_top[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_4[10] = (arbiter_2_4_top[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_3[4] = (arbiter_2_4_top[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_4[1] = (arbiter_2_4_top[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_1[5] = (arbiter_2_4_bottom[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_3[11] = (arbiter_2_4_bottom[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_1_4[8] = (arbiter_2_4_bottom[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_3[2] = (arbiter_2_4_bottom[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_1[9] = (arbiter_3_1_mid[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_2[6] = (arbiter_3_1_mid[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_4[12] = (arbiter_3_1_mid[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_1[0] = (arbiter_3_1_mid[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_4[3] = (arbiter_3_1_mid[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_1[10] = (arbiter_3_1_top[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_2[7] = (arbiter_3_1_top[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_4[13] = (arbiter_3_1_top[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_1[1] = (arbiter_3_1_top[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_4[4] = (arbiter_3_1_top[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_1[8] = (arbiter_3_1_bottom[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_2[5] = (arbiter_3_1_bottom[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_4[11] = (arbiter_3_1_bottom[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_4[2] = (arbiter_3_1_bottom[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_1[12] = (arbiter_3_2_mid[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_2[9] = (arbiter_3_2_mid[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_3[6] = (arbiter_3_2_mid[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_1[3] = (arbiter_3_2_mid[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_2[0] = (arbiter_3_2_mid[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_1[13] = (arbiter_3_2_top[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_2[10] = (arbiter_3_2_top[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_3[7] = (arbiter_3_2_top[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_1[4] = (arbiter_3_2_top[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_2[1] = (arbiter_3_2_top[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_1[11] = (arbiter_3_2_bottom[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_2[8] = (arbiter_3_2_bottom[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_3[5] = (arbiter_3_2_bottom[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_1[2] = (arbiter_3_2_bottom[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_2[12] = (arbiter_3_3_mid[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_3[9] = (arbiter_3_3_mid[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_4[6] = (arbiter_3_3_mid[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_2[3] = (arbiter_3_3_mid[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_3[0] = (arbiter_3_3_mid[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_2[13] = (arbiter_3_3_top[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_3[10] = (arbiter_3_3_top[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_4[7] = (arbiter_3_3_top[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_2[4] = (arbiter_3_3_top[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_3[1] = (arbiter_3_3_top[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_2[11] = (arbiter_3_3_bottom[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_3[8] = (arbiter_3_3_bottom[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_4[5] = (arbiter_3_3_bottom[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_2[2] = (arbiter_3_3_bottom[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_1[6] = (arbiter_3_4_mid[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_3[12] = (arbiter_3_4_mid[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_4[9] = (arbiter_3_4_mid[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_3[3] = (arbiter_3_4_mid[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_4[0] = (arbiter_3_4_mid[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_1[7] = (arbiter_3_4_top[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_3[13] = (arbiter_3_4_top[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_4[10] = (arbiter_3_4_top[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_3[4] = (arbiter_3_4_top[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_4[1] = (arbiter_3_4_top[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_1[5] = (arbiter_3_4_bottom[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_3[11] = (arbiter_3_4_bottom[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_2_4[8] = (arbiter_3_4_bottom[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_3[2] = (arbiter_3_4_bottom[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_1[9] = (arbiter_4_1_mid[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_2[6] = (arbiter_4_1_mid[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_4[12] = (arbiter_4_1_mid[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_1[0] = (arbiter_4_1_mid[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_4[3] = (arbiter_4_1_mid[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_1[10] = (arbiter_4_1_top[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_2[7] = (arbiter_4_1_top[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_4[13] = (arbiter_4_1_top[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_1[1] = (arbiter_4_1_top[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_4[4] = (arbiter_4_1_top[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_1[8] = (arbiter_4_1_bottom[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_2[5] = (arbiter_4_1_bottom[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_4[11] = (arbiter_4_1_bottom[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_4[2] = (arbiter_4_1_bottom[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_1[12] = (arbiter_4_2_mid[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_2[9] = (arbiter_4_2_mid[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_3[6] = (arbiter_4_2_mid[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_1[3] = (arbiter_4_2_mid[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_2[0] = (arbiter_4_2_mid[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_1[13] = (arbiter_4_2_top[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_2[10] = (arbiter_4_2_top[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_3[7] = (arbiter_4_2_top[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_1[4] = (arbiter_4_2_top[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_2[1] = (arbiter_4_2_top[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_1[11] = (arbiter_4_2_bottom[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_2[8] = (arbiter_4_2_bottom[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_3[5] = (arbiter_4_2_bottom[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_1[2] = (arbiter_4_2_bottom[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_2[12] = (arbiter_4_3_mid[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_3[9] = (arbiter_4_3_mid[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_4[6] = (arbiter_4_3_mid[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_2[3] = (arbiter_4_3_mid[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_3[0] = (arbiter_4_3_mid[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_2[13] = (arbiter_4_3_top[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_3[10] = (arbiter_4_3_top[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_4[7] = (arbiter_4_3_top[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_2[4] = (arbiter_4_3_top[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_3[1] = (arbiter_4_3_top[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_2[11] = (arbiter_4_3_bottom[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_3[8] = (arbiter_4_3_bottom[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_4[5] = (arbiter_4_3_bottom[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_2[2] = (arbiter_4_3_bottom[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_1[6] = (arbiter_4_4_mid[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_3[12] = (arbiter_4_4_mid[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_4[9] = (arbiter_4_4_mid[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_3[3] = (arbiter_4_4_mid[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_4[0] = (arbiter_4_4_mid[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_1[7] = (arbiter_4_4_top[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_3[13] = (arbiter_4_4_top[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_4[10] = (arbiter_4_4_top[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_3[4] = (arbiter_4_4_top[3]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_4[1] = (arbiter_4_4_top[4]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_1[5] = (arbiter_4_4_bottom[0]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_3[11] = (arbiter_4_4_bottom[1]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_3_4[8] = (arbiter_4_4_bottom[2]) ? 1'b1 : 1'b0;
	reg_Cell_to_FSM_read_success_bit_4_3[2] = (arbiter_4_4_bottom[3]) ? 1'b1 : 1'b0;
	end

	
	
Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_1_1_mid
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_1_1[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_1_1[0]),
	.addr2(FSM_to_Cell_read_addr_1_4[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_1_4[3]),
	.addr3(FSM_to_Cell_read_addr_4_1[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_4_1[9]),
	.addr4(FSM_to_Cell_read_addr_4_2[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_4_2[6]),
	.addr5(FSM_to_Cell_read_addr_4_4[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_4_4[12]),
	.Arbitration_Result(arbiter_1_1_mid)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_1_1_top
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_1_1[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_1_1[1]),
	.addr2(FSM_to_Cell_read_addr_1_4[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_1_4[4]),
	.addr3(FSM_to_Cell_read_addr_4_1[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_4_1[10]),
	.addr4(FSM_to_Cell_read_addr_4_2[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_4_2[7]),
	.addr5(FSM_to_Cell_read_addr_4_4[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_4_4[13]),
	.Arbitration_Result(arbiter_1_1_top)
);

Read_Addr_Arbiter_Bottom
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_BOTTOM_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_1_1_bottom
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_1_4[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_1_4[2]),
	.addr2(FSM_to_Cell_read_addr_4_1[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_4_1[8]),
	.addr3(FSM_to_Cell_read_addr_4_2[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_4_2[5]),
	.addr4(FSM_to_Cell_read_addr_4_4[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_4_4[11]),
	.Arbitration_Result(arbiter_1_1_bottom)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_1_2_mid
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_1_1[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_1_1[3]),
	.addr2(FSM_to_Cell_read_addr_1_2[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_1_2[0]),
	.addr3(FSM_to_Cell_read_addr_4_1[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_4_1[12]),
	.addr4(FSM_to_Cell_read_addr_4_2[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_4_2[9]),
	.addr5(FSM_to_Cell_read_addr_4_3[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_4_3[6]),
	.Arbitration_Result(arbiter_1_2_mid)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_1_2_top
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_1_1[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_1_1[4]),
	.addr2(FSM_to_Cell_read_addr_1_2[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_1_2[1]),
	.addr3(FSM_to_Cell_read_addr_4_1[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_4_1[13]),
	.addr4(FSM_to_Cell_read_addr_4_2[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_4_2[10]),
	.addr5(FSM_to_Cell_read_addr_4_3[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_4_3[7]),
	.Arbitration_Result(arbiter_1_2_top)
);

Read_Addr_Arbiter_Bottom
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_BOTTOM_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_1_2_bottom
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_1_1[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_1_1[2]),
	.addr2(FSM_to_Cell_read_addr_4_1[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_4_1[11]),
	.addr3(FSM_to_Cell_read_addr_4_2[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_4_2[8]),
	.addr4(FSM_to_Cell_read_addr_4_3[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_4_3[5]),
	.Arbitration_Result(arbiter_1_2_bottom)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_1_3_mid
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_1_2[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_1_2[3]),
	.addr2(FSM_to_Cell_read_addr_1_3[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_1_3[0]),
	.addr3(FSM_to_Cell_read_addr_4_2[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_4_2[12]),
	.addr4(FSM_to_Cell_read_addr_4_3[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_4_3[9]),
	.addr5(FSM_to_Cell_read_addr_4_4[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_4_4[6]),
	.Arbitration_Result(arbiter_1_3_mid)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_1_3_top
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_1_2[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_1_2[4]),
	.addr2(FSM_to_Cell_read_addr_1_3[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_1_3[1]),
	.addr3(FSM_to_Cell_read_addr_4_2[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_4_2[13]),
	.addr4(FSM_to_Cell_read_addr_4_3[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_4_3[10]),
	.addr5(FSM_to_Cell_read_addr_4_4[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_4_4[7]),
	.Arbitration_Result(arbiter_1_3_top)
);

Read_Addr_Arbiter_Bottom
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_BOTTOM_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_1_3_bottom
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_1_2[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_1_2[2]),
	.addr2(FSM_to_Cell_read_addr_4_2[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_4_2[11]),
	.addr3(FSM_to_Cell_read_addr_4_3[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_4_3[8]),
	.addr4(FSM_to_Cell_read_addr_4_4[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_4_4[5]),
	.Arbitration_Result(arbiter_1_3_bottom)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_1_4_mid
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_1_3[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_1_3[3]),
	.addr2(FSM_to_Cell_read_addr_1_4[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_1_4[0]),
	.addr3(FSM_to_Cell_read_addr_4_1[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_4_1[6]),
	.addr4(FSM_to_Cell_read_addr_4_3[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_4_3[12]),
	.addr5(FSM_to_Cell_read_addr_4_4[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_4_4[9]),
	.Arbitration_Result(arbiter_1_4_mid)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_1_4_top
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_1_3[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_1_3[4]),
	.addr2(FSM_to_Cell_read_addr_1_4[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_1_4[1]),
	.addr3(FSM_to_Cell_read_addr_4_1[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_4_1[7]),
	.addr4(FSM_to_Cell_read_addr_4_3[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_4_3[13]),
	.addr5(FSM_to_Cell_read_addr_4_4[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_4_4[10]),
	.Arbitration_Result(arbiter_1_4_top)
);

Read_Addr_Arbiter_Bottom
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_BOTTOM_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_1_4_bottom
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_1_3[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_1_3[2]),
	.addr2(FSM_to_Cell_read_addr_4_1[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_4_1[5]),
	.addr3(FSM_to_Cell_read_addr_4_3[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_4_3[11]),
	.addr4(FSM_to_Cell_read_addr_4_4[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_4_4[8]),
	.Arbitration_Result(arbiter_1_4_bottom)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_2_1_mid
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_1_1[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_1_1[9]),
	.addr2(FSM_to_Cell_read_addr_1_2[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_1_2[6]),
	.addr3(FSM_to_Cell_read_addr_1_4[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_1_4[12]),
	.addr4(FSM_to_Cell_read_addr_2_1[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_2_1[0]),
	.addr5(FSM_to_Cell_read_addr_2_4[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_2_4[3]),
	.Arbitration_Result(arbiter_2_1_mid)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_2_1_top
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_1_1[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_1_1[10]),
	.addr2(FSM_to_Cell_read_addr_1_2[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_1_2[7]),
	.addr3(FSM_to_Cell_read_addr_1_4[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_1_4[13]),
	.addr4(FSM_to_Cell_read_addr_2_1[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_2_1[1]),
	.addr5(FSM_to_Cell_read_addr_2_4[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_2_4[4]),
	.Arbitration_Result(arbiter_2_1_top)
);

Read_Addr_Arbiter_Bottom
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_BOTTOM_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_2_1_bottom
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_1_1[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_1_1[8]),
	.addr2(FSM_to_Cell_read_addr_1_2[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_1_2[5]),
	.addr3(FSM_to_Cell_read_addr_1_4[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_1_4[11]),
	.addr4(FSM_to_Cell_read_addr_2_4[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_2_4[2]),
	.Arbitration_Result(arbiter_2_1_bottom)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_2_2_mid
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_1_1[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_1_1[12]),
	.addr2(FSM_to_Cell_read_addr_1_2[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_1_2[9]),
	.addr3(FSM_to_Cell_read_addr_1_3[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_1_3[6]),
	.addr4(FSM_to_Cell_read_addr_2_1[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_2_1[3]),
	.addr5(FSM_to_Cell_read_addr_2_2[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_2_2[0]),
	.Arbitration_Result(arbiter_2_2_mid)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_2_2_top
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_1_1[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_1_1[13]),
	.addr2(FSM_to_Cell_read_addr_1_2[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_1_2[10]),
	.addr3(FSM_to_Cell_read_addr_1_3[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_1_3[7]),
	.addr4(FSM_to_Cell_read_addr_2_1[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_2_1[4]),
	.addr5(FSM_to_Cell_read_addr_2_2[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_2_2[1]),
	.Arbitration_Result(arbiter_2_2_top)
);

Read_Addr_Arbiter_Bottom
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_BOTTOM_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_2_2_bottom
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_1_1[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_1_1[11]),
	.addr2(FSM_to_Cell_read_addr_1_2[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_1_2[8]),
	.addr3(FSM_to_Cell_read_addr_1_3[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_1_3[5]),
	.addr4(FSM_to_Cell_read_addr_2_1[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_2_1[2]),
	.Arbitration_Result(arbiter_2_2_bottom)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_2_3_mid
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_1_2[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_1_2[12]),
	.addr2(FSM_to_Cell_read_addr_1_3[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_1_3[9]),
	.addr3(FSM_to_Cell_read_addr_1_4[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_1_4[6]),
	.addr4(FSM_to_Cell_read_addr_2_2[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_2_2[3]),
	.addr5(FSM_to_Cell_read_addr_2_3[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_2_3[0]),
	.Arbitration_Result(arbiter_2_3_mid)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_2_3_top
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_1_2[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_1_2[13]),
	.addr2(FSM_to_Cell_read_addr_1_3[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_1_3[10]),
	.addr3(FSM_to_Cell_read_addr_1_4[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_1_4[7]),
	.addr4(FSM_to_Cell_read_addr_2_2[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_2_2[4]),
	.addr5(FSM_to_Cell_read_addr_2_3[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_2_3[1]),
	.Arbitration_Result(arbiter_2_3_top)
);

Read_Addr_Arbiter_Bottom
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_BOTTOM_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_2_3_bottom
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_1_2[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_1_2[11]),
	.addr2(FSM_to_Cell_read_addr_1_3[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_1_3[8]),
	.addr3(FSM_to_Cell_read_addr_1_4[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_1_4[5]),
	.addr4(FSM_to_Cell_read_addr_2_2[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_2_2[2]),
	.Arbitration_Result(arbiter_2_3_bottom)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_2_4_mid
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_1_1[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_1_1[6]),
	.addr2(FSM_to_Cell_read_addr_1_3[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_1_3[12]),
	.addr3(FSM_to_Cell_read_addr_1_4[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_1_4[9]),
	.addr4(FSM_to_Cell_read_addr_2_3[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_2_3[3]),
	.addr5(FSM_to_Cell_read_addr_2_4[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_2_4[0]),
	.Arbitration_Result(arbiter_2_4_mid)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_2_4_top
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_1_1[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_1_1[7]),
	.addr2(FSM_to_Cell_read_addr_1_3[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_1_3[13]),
	.addr3(FSM_to_Cell_read_addr_1_4[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_1_4[10]),
	.addr4(FSM_to_Cell_read_addr_2_3[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_2_3[4]),
	.addr5(FSM_to_Cell_read_addr_2_4[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_2_4[1]),
	.Arbitration_Result(arbiter_2_4_top)
);

Read_Addr_Arbiter_Bottom
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_BOTTOM_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_2_4_bottom
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_1_1[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_1_1[5]),
	.addr2(FSM_to_Cell_read_addr_1_3[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_1_3[11]),
	.addr3(FSM_to_Cell_read_addr_1_4[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_1_4[8]),
	.addr4(FSM_to_Cell_read_addr_2_3[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_2_3[2]),
	.Arbitration_Result(arbiter_2_4_bottom)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_3_1_mid
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_2_1[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_2_1[9]),
	.addr2(FSM_to_Cell_read_addr_2_2[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_2_2[6]),
	.addr3(FSM_to_Cell_read_addr_2_4[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_2_4[12]),
	.addr4(FSM_to_Cell_read_addr_3_1[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_3_1[0]),
	.addr5(FSM_to_Cell_read_addr_3_4[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_3_4[3]),
	.Arbitration_Result(arbiter_3_1_mid)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_3_1_top
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_2_1[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_2_1[10]),
	.addr2(FSM_to_Cell_read_addr_2_2[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_2_2[7]),
	.addr3(FSM_to_Cell_read_addr_2_4[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_2_4[13]),
	.addr4(FSM_to_Cell_read_addr_3_1[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_3_1[1]),
	.addr5(FSM_to_Cell_read_addr_3_4[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_3_4[4]),
	.Arbitration_Result(arbiter_3_1_top)
);

Read_Addr_Arbiter_Bottom
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_BOTTOM_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_3_1_bottom
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_2_1[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_2_1[8]),
	.addr2(FSM_to_Cell_read_addr_2_2[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_2_2[5]),
	.addr3(FSM_to_Cell_read_addr_2_4[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_2_4[11]),
	.addr4(FSM_to_Cell_read_addr_3_4[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_3_4[2]),
	.Arbitration_Result(arbiter_3_1_bottom)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_3_2_mid
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_2_1[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_2_1[12]),
	.addr2(FSM_to_Cell_read_addr_2_2[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_2_2[9]),
	.addr3(FSM_to_Cell_read_addr_2_3[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_2_3[6]),
	.addr4(FSM_to_Cell_read_addr_3_1[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_3_1[3]),
	.addr5(FSM_to_Cell_read_addr_3_2[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_3_2[0]),
	.Arbitration_Result(arbiter_3_2_mid)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_3_2_top
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_2_1[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_2_1[13]),
	.addr2(FSM_to_Cell_read_addr_2_2[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_2_2[10]),
	.addr3(FSM_to_Cell_read_addr_2_3[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_2_3[7]),
	.addr4(FSM_to_Cell_read_addr_3_1[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_3_1[4]),
	.addr5(FSM_to_Cell_read_addr_3_2[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_3_2[1]),
	.Arbitration_Result(arbiter_3_2_top)
);

Read_Addr_Arbiter_Bottom
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_BOTTOM_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_3_2_bottom
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_2_1[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_2_1[11]),
	.addr2(FSM_to_Cell_read_addr_2_2[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_2_2[8]),
	.addr3(FSM_to_Cell_read_addr_2_3[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_2_3[5]),
	.addr4(FSM_to_Cell_read_addr_3_1[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_3_1[2]),
	.Arbitration_Result(arbiter_3_2_bottom)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_3_3_mid
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_2_2[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_2_2[12]),
	.addr2(FSM_to_Cell_read_addr_2_3[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_2_3[9]),
	.addr3(FSM_to_Cell_read_addr_2_4[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_2_4[6]),
	.addr4(FSM_to_Cell_read_addr_3_2[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_3_2[3]),
	.addr5(FSM_to_Cell_read_addr_3_3[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_3_3[0]),
	.Arbitration_Result(arbiter_3_3_mid)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_3_3_top
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_2_2[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_2_2[13]),
	.addr2(FSM_to_Cell_read_addr_2_3[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_2_3[10]),
	.addr3(FSM_to_Cell_read_addr_2_4[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_2_4[7]),
	.addr4(FSM_to_Cell_read_addr_3_2[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_3_2[4]),
	.addr5(FSM_to_Cell_read_addr_3_3[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_3_3[1]),
	.Arbitration_Result(arbiter_3_3_top)
);

Read_Addr_Arbiter_Bottom
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_BOTTOM_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_3_3_bottom
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_2_2[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_2_2[11]),
	.addr2(FSM_to_Cell_read_addr_2_3[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_2_3[8]),
	.addr3(FSM_to_Cell_read_addr_2_4[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_2_4[5]),
	.addr4(FSM_to_Cell_read_addr_3_2[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_3_2[2]),
	.Arbitration_Result(arbiter_3_3_bottom)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_3_4_mid
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_2_1[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_2_1[6]),
	.addr2(FSM_to_Cell_read_addr_2_3[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_2_3[12]),
	.addr3(FSM_to_Cell_read_addr_2_4[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_2_4[9]),
	.addr4(FSM_to_Cell_read_addr_3_3[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_3_3[3]),
	.addr5(FSM_to_Cell_read_addr_3_4[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_3_4[0]),
	.Arbitration_Result(arbiter_3_4_mid)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_3_4_top
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_2_1[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_2_1[7]),
	.addr2(FSM_to_Cell_read_addr_2_3[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_2_3[13]),
	.addr3(FSM_to_Cell_read_addr_2_4[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_2_4[10]),
	.addr4(FSM_to_Cell_read_addr_3_3[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_3_3[4]),
	.addr5(FSM_to_Cell_read_addr_3_4[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_3_4[1]),
	.Arbitration_Result(arbiter_3_4_top)
);

Read_Addr_Arbiter_Bottom
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_BOTTOM_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_3_4_bottom
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_2_1[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_2_1[5]),
	.addr2(FSM_to_Cell_read_addr_2_3[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_2_3[11]),
	.addr3(FSM_to_Cell_read_addr_2_4[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_2_4[8]),
	.addr4(FSM_to_Cell_read_addr_3_3[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_3_3[2]),
	.Arbitration_Result(arbiter_3_4_bottom)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_4_1_mid
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_3_1[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_3_1[9]),
	.addr2(FSM_to_Cell_read_addr_3_2[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_3_2[6]),
	.addr3(FSM_to_Cell_read_addr_3_4[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_3_4[12]),
	.addr4(FSM_to_Cell_read_addr_4_1[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_4_1[0]),
	.addr5(FSM_to_Cell_read_addr_4_4[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_4_4[3]),
	.Arbitration_Result(arbiter_4_1_mid)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_4_1_top
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_3_1[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_3_1[10]),
	.addr2(FSM_to_Cell_read_addr_3_2[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_3_2[7]),
	.addr3(FSM_to_Cell_read_addr_3_4[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_3_4[13]),
	.addr4(FSM_to_Cell_read_addr_4_1[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_4_1[1]),
	.addr5(FSM_to_Cell_read_addr_4_4[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_4_4[4]),
	.Arbitration_Result(arbiter_4_1_top)
);

Read_Addr_Arbiter_Bottom
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_BOTTOM_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_4_1_bottom
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_3_1[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_3_1[8]),
	.addr2(FSM_to_Cell_read_addr_3_2[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_3_2[5]),
	.addr3(FSM_to_Cell_read_addr_3_4[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_3_4[11]),
	.addr4(FSM_to_Cell_read_addr_4_4[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_4_4[2]),
	.Arbitration_Result(arbiter_4_1_bottom)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_4_2_mid
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_3_1[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_3_1[12]),
	.addr2(FSM_to_Cell_read_addr_3_2[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_3_2[9]),
	.addr3(FSM_to_Cell_read_addr_3_3[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_3_3[6]),
	.addr4(FSM_to_Cell_read_addr_4_1[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_4_1[3]),
	.addr5(FSM_to_Cell_read_addr_4_2[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_4_2[0]),
	.Arbitration_Result(arbiter_4_2_mid)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_4_2_top
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_3_1[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_3_1[13]),
	.addr2(FSM_to_Cell_read_addr_3_2[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_3_2[10]),
	.addr3(FSM_to_Cell_read_addr_3_3[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_3_3[7]),
	.addr4(FSM_to_Cell_read_addr_4_1[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_4_1[4]),
	.addr5(FSM_to_Cell_read_addr_4_2[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_4_2[1]),
	.Arbitration_Result(arbiter_4_2_top)
);

Read_Addr_Arbiter_Bottom
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_BOTTOM_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_4_2_bottom
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_3_1[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_3_1[11]),
	.addr2(FSM_to_Cell_read_addr_3_2[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_3_2[8]),
	.addr3(FSM_to_Cell_read_addr_3_3[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_3_3[5]),
	.addr4(FSM_to_Cell_read_addr_4_1[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_4_1[2]),
	.Arbitration_Result(arbiter_4_2_bottom)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_4_3_mid
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_3_2[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_3_2[12]),
	.addr2(FSM_to_Cell_read_addr_3_3[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_3_3[9]),
	.addr3(FSM_to_Cell_read_addr_3_4[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_3_4[6]),
	.addr4(FSM_to_Cell_read_addr_4_2[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_4_2[3]),
	.addr5(FSM_to_Cell_read_addr_4_3[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_4_3[0]),
	.Arbitration_Result(arbiter_4_3_mid)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_4_3_top
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_3_2[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_3_2[13]),
	.addr2(FSM_to_Cell_read_addr_3_3[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_3_3[10]),
	.addr3(FSM_to_Cell_read_addr_3_4[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_3_4[7]),
	.addr4(FSM_to_Cell_read_addr_4_2[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_4_2[4]),
	.addr5(FSM_to_Cell_read_addr_4_3[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_4_3[1]),
	.Arbitration_Result(arbiter_4_3_top)
);

Read_Addr_Arbiter_Bottom
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_BOTTOM_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_4_3_bottom
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_3_2[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_3_2[11]),
	.addr2(FSM_to_Cell_read_addr_3_3[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_3_3[8]),
	.addr3(FSM_to_Cell_read_addr_3_4[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_3_4[5]),
	.addr4(FSM_to_Cell_read_addr_4_2[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_4_2[2]),
	.Arbitration_Result(arbiter_4_3_bottom)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_4_4_mid
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_3_1[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_3_1[6]),
	.addr2(FSM_to_Cell_read_addr_3_3[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_3_3[12]),
	.addr3(FSM_to_Cell_read_addr_3_4[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_3_4[9]),
	.addr4(FSM_to_Cell_read_addr_4_3[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_4_3[3]),
	.addr5(FSM_to_Cell_read_addr_4_4[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_4_4[0]),
	.Arbitration_Result(arbiter_4_4_mid)
);

Read_Addr_Arbiter
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_4_4_top
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_3_1[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_3_1[7]),
	.addr2(FSM_to_Cell_read_addr_3_3[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_3_3[13]),
	.addr3(FSM_to_Cell_read_addr_3_4[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_3_4[10]),
	.addr4(FSM_to_Cell_read_addr_4_3[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_4_3[4]),
	.addr5(FSM_to_Cell_read_addr_4_4[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH]),
	.enable5(enable_reading_4_4[1]),
	.Arbitration_Result(arbiter_4_4_top)
);

Read_Addr_Arbiter_Bottom
#(
	.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),
	.RDADDR_ARBITER_SIZE(RDADDR_ARBITER_BOTTOM_SIZE),
	.RDADDR_ARBITER_MSB(RDADDR_ARBITER_MSB)
)
Read_Addr_Arbiter_4_4_bottom
(
	.clk(clk),
	.rst(rst),
	.addr1(FSM_to_Cell_read_addr_3_1[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH]),
	.enable1(enable_reading_3_1[5]),
	.addr2(FSM_to_Cell_read_addr_3_3[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH]),
	.enable2(enable_reading_3_3[11]),
	.addr3(FSM_to_Cell_read_addr_3_4[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH]),
	.enable3(enable_reading_3_4[8]),
	.addr4(FSM_to_Cell_read_addr_4_3[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH]),
	.enable4(enable_reading_4_3[2]),
	.Arbitration_Result(arbiter_4_4_bottom)
);


endmodule