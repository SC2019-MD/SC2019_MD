/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Module: fp_mult.v
//
//	Function:
//				Wrapper on top of FP_MUL, to meet the port configuration in the old design
//
// Dependency:
//				FP_MUL.v
//
// Latency: 4 cycles

//
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module fp_mult
#(
	parameter DATA_WIDTH = 32
)
(
	input clk,
	input [DATA_WIDTH-1:0] in1,
	input [DATA_WIDTH-1:0] in2,
	output [DATA_WIDTH-1:0] result
);

	FP_MUL FP_MUL
	(
		.clk(clk),
		.ena(1'b1),
		.clr(1'b0),
		.ay(in1),
		.az(in2),
		.result(result)
	);

endmodule
