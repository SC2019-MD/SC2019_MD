module Pipeline_local_to_global_mapping
#(
	parameter DATA_WIDTH							= 32,
	parameter NUM_NEIGHBOR_CELLS				= 13,
	parameter TOTAL_CELL_NUM					= 64,
	parameter CELL_ADDR_WIDTH					= 7,
	parameter CELL_ID_WIDTH						= 3,
	parameter PARTICLE_ID_WIDTH				= CELL_ID_WIDTH*3+CELL_ADDR_WIDTH
)
(
	input clk, 
	input rst, 
	input [TOTAL_CELL_NUM*3*DATA_WIDTH-1:0] Position_Cache_readout_position,
	input [(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:0] FSM_to_Cell_read_addr_1_1,
	input FSM_to_Cell_rden_1_1,
	input [CELL_ID_WIDTH-1:0] cellz_1_1,
	
	// Force cache mapping
	input [PARTICLE_ID_WIDTH-1:0] ref_particle_id_1_1,
	input [DATA_WIDTH-1:0] ref_LJ_Force_X_1_1,
	input [DATA_WIDTH-1:0] ref_LJ_Force_Y_1_1,
	input [DATA_WIDTH-1:0] ref_LJ_Force_Z_1_1,
	input ref_forceoutput_valid_1_1,
	input [PARTICLE_ID_WIDTH-1:0] neighbor_particle_id_1_1,
	input [DATA_WIDTH-1:0] neighbor_LJ_Force_X_1_1,
	input [DATA_WIDTH-1:0] neighbor_LJ_Force_Y_1_1,
	input [DATA_WIDTH-1:0] neighbor_LJ_Force_Z_1_1,
	input neighbor_forceoutput_valid_1_1,
	
	
	output [(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH-1:0] cells_to_pipeline_1_1,
	output [TOTAL_CELL_NUM*CELL_ADDR_WIDTH-1:0] FSM_to_Cell_read_addr,
	output [TOTAL_CELL_NUM-1:0] FSM_to_Cell_rden,
	
	// Force cache mapping
	output [TOTAL_CELL_NUM-1:0] to_force_cache_partial_force_valid,
	output [TOTAL_CELL_NUM*PARTICLE_ID_WIDTH-1:0] to_force_cache_particle_id,
	output [TOTAL_CELL_NUM*DATA_WIDTH-1:0] to_force_cache_LJ_Force_Z,
	output [TOTAL_CELL_NUM*DATA_WIDTH-1:0] to_force_cache_LJ_Force_Y,
	output [TOTAL_CELL_NUM*DATA_WIDTH-1:0] to_force_cache_LJ_Force_X
);

reg [(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH-1:0] reg_cells_to_pipeline_1_1;
reg [TOTAL_CELL_NUM*CELL_ADDR_WIDTH-1:0] reg_FSM_to_Cell_read_addr;
reg [TOTAL_CELL_NUM-1:0] reg_FSM_to_Cell_rden;
reg [TOTAL_CELL_NUM-1:0] reg_to_force_cache_partial_force_valid;
reg [TOTAL_CELL_NUM*PARTICLE_ID_WIDTH-1:0] reg_to_force_cache_particle_id;
reg [TOTAL_CELL_NUM*DATA_WIDTH-1:0] reg_to_force_cache_LJ_Force_Z;
reg [TOTAL_CELL_NUM*DATA_WIDTH-1:0] reg_to_force_cache_LJ_Force_Y;
reg [TOTAL_CELL_NUM*DATA_WIDTH-1:0] reg_to_force_cache_LJ_Force_X;
assign cells_to_pipeline_1_1 = reg_cells_to_pipeline_1_1;
assign FSM_to_Cell_read_addr = reg_FSM_to_Cell_read_addr;
assign FSM_to_Cell_rden = reg_FSM_to_Cell_rden;
assign to_force_cache_partial_force_valid = reg_to_force_cache_partial_force_valid;
assign to_force_cache_particle_id = reg_to_force_cache_particle_id;
assign to_force_cache_LJ_Force_Z = reg_to_force_cache_LJ_Force_Z;
assign to_force_cache_LJ_Force_Y = reg_to_force_cache_LJ_Force_Y;
assign to_force_cache_LJ_Force_X = reg_to_force_cache_LJ_Force_X;


always@(*)
	begin
	if (rst)
		begin
		reg_cells_to_pipeline_1_1 <= 0;
		reg_FSM_to_Cell_read_addr <= 0;
		reg_FSM_to_Cell_rden <= 0;
		reg_to_force_cache_partial_force_valid <= 0;
		reg_to_force_cache_particle_id <= 0;
		reg_to_force_cache_LJ_Force_Z <= 0;
		reg_to_force_cache_LJ_Force_Y <= 0;
		reg_to_force_cache_LJ_Force_X <= 0;
		end
	else
		begin
		case(cellz_1_1)
			1:
				begin
				reg_to_force_cache_LJ_Force_Z[1*DATA_WIDTH-1:0*DATA_WIDTH] <= ref_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[2*DATA_WIDTH-1:1*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[3*DATA_WIDTH-1:2*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[4*DATA_WIDTH-1:3*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[5*DATA_WIDTH-1:4*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[6*DATA_WIDTH-1:5*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[7*DATA_WIDTH-1:6*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[8*DATA_WIDTH-1:7*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[9*DATA_WIDTH-1:8*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[10*DATA_WIDTH-1:9*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[11*DATA_WIDTH-1:10*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[12*DATA_WIDTH-1:11*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[13*DATA_WIDTH-1:12*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[14*DATA_WIDTH-1:13*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[15*DATA_WIDTH-1:14*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[16*DATA_WIDTH-1:15*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[17*DATA_WIDTH-1:16*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[18*DATA_WIDTH-1:17*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[19*DATA_WIDTH-1:18*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[20*DATA_WIDTH-1:19*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[21*DATA_WIDTH-1:20*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[22*DATA_WIDTH-1:21*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[23*DATA_WIDTH-1:22*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[24*DATA_WIDTH-1:23*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[25*DATA_WIDTH-1:24*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[26*DATA_WIDTH-1:25*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[27*DATA_WIDTH-1:26*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[28*DATA_WIDTH-1:27*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[29*DATA_WIDTH-1:28*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[30*DATA_WIDTH-1:29*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[31*DATA_WIDTH-1:30*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[32*DATA_WIDTH-1:31*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[33*DATA_WIDTH-1:32*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[34*DATA_WIDTH-1:33*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[35*DATA_WIDTH-1:34*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[36*DATA_WIDTH-1:35*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[37*DATA_WIDTH-1:36*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[38*DATA_WIDTH-1:37*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[39*DATA_WIDTH-1:38*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[40*DATA_WIDTH-1:39*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[41*DATA_WIDTH-1:40*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[42*DATA_WIDTH-1:41*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[43*DATA_WIDTH-1:42*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[44*DATA_WIDTH-1:43*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[45*DATA_WIDTH-1:44*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[46*DATA_WIDTH-1:45*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[47*DATA_WIDTH-1:46*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[48*DATA_WIDTH-1:47*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[49*DATA_WIDTH-1:48*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[50*DATA_WIDTH-1:49*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[51*DATA_WIDTH-1:50*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[52*DATA_WIDTH-1:51*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[53*DATA_WIDTH-1:52*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[54*DATA_WIDTH-1:53*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[55*DATA_WIDTH-1:54*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[56*DATA_WIDTH-1:55*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[57*DATA_WIDTH-1:56*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[58*DATA_WIDTH-1:57*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[59*DATA_WIDTH-1:58*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[60*DATA_WIDTH-1:59*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[61*DATA_WIDTH-1:60*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[62*DATA_WIDTH-1:61*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[63*DATA_WIDTH-1:62*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[64*DATA_WIDTH-1:63*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[1*DATA_WIDTH-1:0*DATA_WIDTH] <= ref_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[2*DATA_WIDTH-1:1*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[3*DATA_WIDTH-1:2*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[4*DATA_WIDTH-1:3*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[5*DATA_WIDTH-1:4*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[6*DATA_WIDTH-1:5*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[7*DATA_WIDTH-1:6*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[8*DATA_WIDTH-1:7*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[9*DATA_WIDTH-1:8*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[10*DATA_WIDTH-1:9*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[11*DATA_WIDTH-1:10*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[12*DATA_WIDTH-1:11*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[13*DATA_WIDTH-1:12*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[14*DATA_WIDTH-1:13*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[15*DATA_WIDTH-1:14*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[16*DATA_WIDTH-1:15*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[17*DATA_WIDTH-1:16*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[18*DATA_WIDTH-1:17*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[19*DATA_WIDTH-1:18*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[20*DATA_WIDTH-1:19*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[21*DATA_WIDTH-1:20*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[22*DATA_WIDTH-1:21*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[23*DATA_WIDTH-1:22*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[24*DATA_WIDTH-1:23*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[25*DATA_WIDTH-1:24*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[26*DATA_WIDTH-1:25*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[27*DATA_WIDTH-1:26*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[28*DATA_WIDTH-1:27*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[29*DATA_WIDTH-1:28*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[30*DATA_WIDTH-1:29*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[31*DATA_WIDTH-1:30*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[32*DATA_WIDTH-1:31*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[33*DATA_WIDTH-1:32*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[34*DATA_WIDTH-1:33*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[35*DATA_WIDTH-1:34*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[36*DATA_WIDTH-1:35*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[37*DATA_WIDTH-1:36*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[38*DATA_WIDTH-1:37*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[39*DATA_WIDTH-1:38*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[40*DATA_WIDTH-1:39*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[41*DATA_WIDTH-1:40*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[42*DATA_WIDTH-1:41*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[43*DATA_WIDTH-1:42*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[44*DATA_WIDTH-1:43*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[45*DATA_WIDTH-1:44*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[46*DATA_WIDTH-1:45*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[47*DATA_WIDTH-1:46*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[48*DATA_WIDTH-1:47*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[49*DATA_WIDTH-1:48*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[50*DATA_WIDTH-1:49*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[51*DATA_WIDTH-1:50*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[52*DATA_WIDTH-1:51*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[53*DATA_WIDTH-1:52*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[54*DATA_WIDTH-1:53*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[55*DATA_WIDTH-1:54*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[56*DATA_WIDTH-1:55*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[57*DATA_WIDTH-1:56*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[58*DATA_WIDTH-1:57*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[59*DATA_WIDTH-1:58*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[60*DATA_WIDTH-1:59*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[61*DATA_WIDTH-1:60*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[62*DATA_WIDTH-1:61*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[63*DATA_WIDTH-1:62*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[64*DATA_WIDTH-1:63*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[1*DATA_WIDTH-1:0*DATA_WIDTH] <= ref_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[2*DATA_WIDTH-1:1*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[3*DATA_WIDTH-1:2*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[4*DATA_WIDTH-1:3*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[5*DATA_WIDTH-1:4*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[6*DATA_WIDTH-1:5*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[7*DATA_WIDTH-1:6*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[8*DATA_WIDTH-1:7*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[9*DATA_WIDTH-1:8*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[10*DATA_WIDTH-1:9*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[11*DATA_WIDTH-1:10*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[12*DATA_WIDTH-1:11*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[13*DATA_WIDTH-1:12*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[14*DATA_WIDTH-1:13*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[15*DATA_WIDTH-1:14*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[16*DATA_WIDTH-1:15*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[17*DATA_WIDTH-1:16*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[18*DATA_WIDTH-1:17*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[19*DATA_WIDTH-1:18*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[20*DATA_WIDTH-1:19*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[21*DATA_WIDTH-1:20*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[22*DATA_WIDTH-1:21*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[23*DATA_WIDTH-1:22*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[24*DATA_WIDTH-1:23*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[25*DATA_WIDTH-1:24*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[26*DATA_WIDTH-1:25*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[27*DATA_WIDTH-1:26*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[28*DATA_WIDTH-1:27*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[29*DATA_WIDTH-1:28*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[30*DATA_WIDTH-1:29*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[31*DATA_WIDTH-1:30*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[32*DATA_WIDTH-1:31*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[33*DATA_WIDTH-1:32*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[34*DATA_WIDTH-1:33*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[35*DATA_WIDTH-1:34*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[36*DATA_WIDTH-1:35*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[37*DATA_WIDTH-1:36*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[38*DATA_WIDTH-1:37*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[39*DATA_WIDTH-1:38*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[40*DATA_WIDTH-1:39*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[41*DATA_WIDTH-1:40*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[42*DATA_WIDTH-1:41*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[43*DATA_WIDTH-1:42*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[44*DATA_WIDTH-1:43*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[45*DATA_WIDTH-1:44*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[46*DATA_WIDTH-1:45*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[47*DATA_WIDTH-1:46*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[48*DATA_WIDTH-1:47*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[49*DATA_WIDTH-1:48*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[50*DATA_WIDTH-1:49*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[51*DATA_WIDTH-1:50*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[52*DATA_WIDTH-1:51*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[53*DATA_WIDTH-1:52*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[54*DATA_WIDTH-1:53*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[55*DATA_WIDTH-1:54*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[56*DATA_WIDTH-1:55*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[57*DATA_WIDTH-1:56*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[58*DATA_WIDTH-1:57*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[59*DATA_WIDTH-1:58*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[60*DATA_WIDTH-1:59*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[61*DATA_WIDTH-1:60*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[62*DATA_WIDTH-1:61*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[63*DATA_WIDTH-1:62*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[64*DATA_WIDTH-1:63*DATA_WIDTH] <= 0;
				reg_to_force_cache_particle_id[1*PARTICLE_ID_WIDTH-1:0*PARTICLE_ID_WIDTH] <= ref_particle_id_1_1;
				reg_to_force_cache_particle_id[2*PARTICLE_ID_WIDTH-1:1*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[3*PARTICLE_ID_WIDTH-1:2*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[4*PARTICLE_ID_WIDTH-1:3*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[5*PARTICLE_ID_WIDTH-1:4*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[6*PARTICLE_ID_WIDTH-1:5*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[7*PARTICLE_ID_WIDTH-1:6*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[8*PARTICLE_ID_WIDTH-1:7*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[9*PARTICLE_ID_WIDTH-1:8*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[10*PARTICLE_ID_WIDTH-1:9*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[11*PARTICLE_ID_WIDTH-1:10*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[12*PARTICLE_ID_WIDTH-1:11*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[13*PARTICLE_ID_WIDTH-1:12*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[14*PARTICLE_ID_WIDTH-1:13*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[15*PARTICLE_ID_WIDTH-1:14*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[16*PARTICLE_ID_WIDTH-1:15*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[17*PARTICLE_ID_WIDTH-1:16*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[18*PARTICLE_ID_WIDTH-1:17*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[19*PARTICLE_ID_WIDTH-1:18*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[20*PARTICLE_ID_WIDTH-1:19*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[21*PARTICLE_ID_WIDTH-1:20*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[22*PARTICLE_ID_WIDTH-1:21*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[23*PARTICLE_ID_WIDTH-1:22*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[24*PARTICLE_ID_WIDTH-1:23*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[25*PARTICLE_ID_WIDTH-1:24*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[26*PARTICLE_ID_WIDTH-1:25*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[27*PARTICLE_ID_WIDTH-1:26*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[28*PARTICLE_ID_WIDTH-1:27*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[29*PARTICLE_ID_WIDTH-1:28*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[30*PARTICLE_ID_WIDTH-1:29*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[31*PARTICLE_ID_WIDTH-1:30*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[32*PARTICLE_ID_WIDTH-1:31*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[33*PARTICLE_ID_WIDTH-1:32*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[34*PARTICLE_ID_WIDTH-1:33*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[35*PARTICLE_ID_WIDTH-1:34*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[36*PARTICLE_ID_WIDTH-1:35*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[37*PARTICLE_ID_WIDTH-1:36*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[38*PARTICLE_ID_WIDTH-1:37*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[39*PARTICLE_ID_WIDTH-1:38*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[40*PARTICLE_ID_WIDTH-1:39*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[41*PARTICLE_ID_WIDTH-1:40*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[42*PARTICLE_ID_WIDTH-1:41*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[43*PARTICLE_ID_WIDTH-1:42*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[44*PARTICLE_ID_WIDTH-1:43*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[45*PARTICLE_ID_WIDTH-1:44*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[46*PARTICLE_ID_WIDTH-1:45*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[47*PARTICLE_ID_WIDTH-1:46*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[48*PARTICLE_ID_WIDTH-1:47*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[49*PARTICLE_ID_WIDTH-1:48*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[50*PARTICLE_ID_WIDTH-1:49*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[51*PARTICLE_ID_WIDTH-1:50*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[52*PARTICLE_ID_WIDTH-1:51*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[53*PARTICLE_ID_WIDTH-1:52*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[54*PARTICLE_ID_WIDTH-1:53*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[55*PARTICLE_ID_WIDTH-1:54*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[56*PARTICLE_ID_WIDTH-1:55*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[57*PARTICLE_ID_WIDTH-1:56*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[58*PARTICLE_ID_WIDTH-1:57*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[59*PARTICLE_ID_WIDTH-1:58*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[60*PARTICLE_ID_WIDTH-1:59*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[61*PARTICLE_ID_WIDTH-1:60*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[62*PARTICLE_ID_WIDTH-1:61*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[63*PARTICLE_ID_WIDTH-1:62*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[64*PARTICLE_ID_WIDTH-1:63*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_partial_force_valid[0] <= ref_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[1] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[2] <= 1'b0;
				reg_to_force_cache_partial_force_valid[3] <= 1'b0;
				reg_to_force_cache_partial_force_valid[4] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[5] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[6] <= 1'b0;
				reg_to_force_cache_partial_force_valid[7] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[8] <= 1'b0;
				reg_to_force_cache_partial_force_valid[9] <= 1'b0;
				reg_to_force_cache_partial_force_valid[10] <= 1'b0;
				reg_to_force_cache_partial_force_valid[11] <= 1'b0;
				reg_to_force_cache_partial_force_valid[12] <= 1'b0;
				reg_to_force_cache_partial_force_valid[13] <= 1'b0;
				reg_to_force_cache_partial_force_valid[14] <= 1'b0;
				reg_to_force_cache_partial_force_valid[15] <= 1'b0;
				reg_to_force_cache_partial_force_valid[16] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[17] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[18] <= 1'b0;
				reg_to_force_cache_partial_force_valid[19] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[20] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[21] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[22] <= 1'b0;
				reg_to_force_cache_partial_force_valid[23] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[24] <= 1'b0;
				reg_to_force_cache_partial_force_valid[25] <= 1'b0;
				reg_to_force_cache_partial_force_valid[26] <= 1'b0;
				reg_to_force_cache_partial_force_valid[27] <= 1'b0;
				reg_to_force_cache_partial_force_valid[28] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[29] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[30] <= 1'b0;
				reg_to_force_cache_partial_force_valid[31] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[32] <= 1'b0;
				reg_to_force_cache_partial_force_valid[33] <= 1'b0;
				reg_to_force_cache_partial_force_valid[34] <= 1'b0;
				reg_to_force_cache_partial_force_valid[35] <= 1'b0;
				reg_to_force_cache_partial_force_valid[36] <= 1'b0;
				reg_to_force_cache_partial_force_valid[37] <= 1'b0;
				reg_to_force_cache_partial_force_valid[38] <= 1'b0;
				reg_to_force_cache_partial_force_valid[39] <= 1'b0;
				reg_to_force_cache_partial_force_valid[40] <= 1'b0;
				reg_to_force_cache_partial_force_valid[41] <= 1'b0;
				reg_to_force_cache_partial_force_valid[42] <= 1'b0;
				reg_to_force_cache_partial_force_valid[43] <= 1'b0;
				reg_to_force_cache_partial_force_valid[44] <= 1'b0;
				reg_to_force_cache_partial_force_valid[45] <= 1'b0;
				reg_to_force_cache_partial_force_valid[46] <= 1'b0;
				reg_to_force_cache_partial_force_valid[47] <= 1'b0;
				reg_to_force_cache_partial_force_valid[48] <= 1'b0;
				reg_to_force_cache_partial_force_valid[49] <= 1'b0;
				reg_to_force_cache_partial_force_valid[50] <= 1'b0;
				reg_to_force_cache_partial_force_valid[51] <= 1'b0;
				reg_to_force_cache_partial_force_valid[52] <= 1'b0;
				reg_to_force_cache_partial_force_valid[53] <= 1'b0;
				reg_to_force_cache_partial_force_valid[54] <= 1'b0;
				reg_to_force_cache_partial_force_valid[55] <= 1'b0;
				reg_to_force_cache_partial_force_valid[56] <= 1'b0;
				reg_to_force_cache_partial_force_valid[57] <= 1'b0;
				reg_to_force_cache_partial_force_valid[58] <= 1'b0;
				reg_to_force_cache_partial_force_valid[59] <= 1'b0;
				reg_to_force_cache_partial_force_valid[60] <= 1'b0;
				reg_to_force_cache_partial_force_valid[61] <= 1'b0;
				reg_to_force_cache_partial_force_valid[62] <= 1'b0;
				reg_to_force_cache_partial_force_valid[63] <= 1'b0;
				reg_cells_to_pipeline_1_1 <= 	{
														Position_Cache_readout_position[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH],
														Position_Cache_readout_position[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH],
														Position_Cache_readout_position[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH],
														Position_Cache_readout_position[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH],
														Position_Cache_readout_position[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH],
														Position_Cache_readout_position[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH],
														Position_Cache_readout_position[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH],
														Position_Cache_readout_position[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH],
														Position_Cache_readout_position[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH],
														Position_Cache_readout_position[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH],
														Position_Cache_readout_position[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH],
														Position_Cache_readout_position[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH],
														Position_Cache_readout_position[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH],
														Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH]
														};
				reg_FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[15*CELL_ADDR_WIDTH-1:14*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[16*CELL_ADDR_WIDTH-1:15*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[17*CELL_ADDR_WIDTH-1:16*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[18*CELL_ADDR_WIDTH-1:17*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[19*CELL_ADDR_WIDTH-1:18*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[20*CELL_ADDR_WIDTH-1:19*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[21*CELL_ADDR_WIDTH-1:20*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[22*CELL_ADDR_WIDTH-1:21*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[23*CELL_ADDR_WIDTH-1:22*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[24*CELL_ADDR_WIDTH-1:23*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[25*CELL_ADDR_WIDTH-1:24*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[26*CELL_ADDR_WIDTH-1:25*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[27*CELL_ADDR_WIDTH-1:26*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[28*CELL_ADDR_WIDTH-1:27*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[29*CELL_ADDR_WIDTH-1:28*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[30*CELL_ADDR_WIDTH-1:29*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[31*CELL_ADDR_WIDTH-1:30*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[32*CELL_ADDR_WIDTH-1:31*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[33*CELL_ADDR_WIDTH-1:32*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[34*CELL_ADDR_WIDTH-1:33*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[35*CELL_ADDR_WIDTH-1:34*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[36*CELL_ADDR_WIDTH-1:35*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[37*CELL_ADDR_WIDTH-1:36*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[38*CELL_ADDR_WIDTH-1:37*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[39*CELL_ADDR_WIDTH-1:38*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[40*CELL_ADDR_WIDTH-1:39*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[41*CELL_ADDR_WIDTH-1:40*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[42*CELL_ADDR_WIDTH-1:41*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[43*CELL_ADDR_WIDTH-1:42*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[44*CELL_ADDR_WIDTH-1:43*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[45*CELL_ADDR_WIDTH-1:44*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[46*CELL_ADDR_WIDTH-1:45*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[47*CELL_ADDR_WIDTH-1:46*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[48*CELL_ADDR_WIDTH-1:47*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[49*CELL_ADDR_WIDTH-1:48*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[50*CELL_ADDR_WIDTH-1:49*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[51*CELL_ADDR_WIDTH-1:50*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[52*CELL_ADDR_WIDTH-1:51*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[53*CELL_ADDR_WIDTH-1:52*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[54*CELL_ADDR_WIDTH-1:53*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[55*CELL_ADDR_WIDTH-1:54*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[56*CELL_ADDR_WIDTH-1:55*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[57*CELL_ADDR_WIDTH-1:56*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[58*CELL_ADDR_WIDTH-1:57*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[59*CELL_ADDR_WIDTH-1:58*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[60*CELL_ADDR_WIDTH-1:59*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[61*CELL_ADDR_WIDTH-1:60*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[62*CELL_ADDR_WIDTH-1:61*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[63*CELL_ADDR_WIDTH-1:62*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[64*CELL_ADDR_WIDTH-1:63*CELL_ADDR_WIDTH] <= 0;
				if (FSM_to_Cell_rden_1_1)
					begin
					reg_FSM_to_Cell_rden[0] <= 1'b1;
					reg_FSM_to_Cell_rden[1] <= 1'b1;
					reg_FSM_to_Cell_rden[2] <= 1'b0;
					reg_FSM_to_Cell_rden[3] <= 1'b0;
					reg_FSM_to_Cell_rden[4] <= 1'b1;
					reg_FSM_to_Cell_rden[5] <= 1'b1;
					reg_FSM_to_Cell_rden[6] <= 1'b0;
					reg_FSM_to_Cell_rden[7] <= 1'b1;
					reg_FSM_to_Cell_rden[8] <= 1'b0;
					reg_FSM_to_Cell_rden[9] <= 1'b0;
					reg_FSM_to_Cell_rden[10] <= 1'b0;
					reg_FSM_to_Cell_rden[11] <= 1'b0;
					reg_FSM_to_Cell_rden[12] <= 1'b0;
					reg_FSM_to_Cell_rden[13] <= 1'b0;
					reg_FSM_to_Cell_rden[14] <= 1'b0;
					reg_FSM_to_Cell_rden[15] <= 1'b0;
					reg_FSM_to_Cell_rden[16] <= 1'b1;
					reg_FSM_to_Cell_rden[17] <= 1'b1;
					reg_FSM_to_Cell_rden[18] <= 1'b0;
					reg_FSM_to_Cell_rden[19] <= 1'b1;
					reg_FSM_to_Cell_rden[20] <= 1'b1;
					reg_FSM_to_Cell_rden[21] <= 1'b1;
					reg_FSM_to_Cell_rden[22] <= 1'b0;
					reg_FSM_to_Cell_rden[23] <= 1'b1;
					reg_FSM_to_Cell_rden[24] <= 1'b0;
					reg_FSM_to_Cell_rden[25] <= 1'b0;
					reg_FSM_to_Cell_rden[26] <= 1'b0;
					reg_FSM_to_Cell_rden[27] <= 1'b0;
					reg_FSM_to_Cell_rden[28] <= 1'b1;
					reg_FSM_to_Cell_rden[29] <= 1'b1;
					reg_FSM_to_Cell_rden[30] <= 1'b0;
					reg_FSM_to_Cell_rden[31] <= 1'b1;
					reg_FSM_to_Cell_rden[32] <= 1'b0;
					reg_FSM_to_Cell_rden[33] <= 1'b0;
					reg_FSM_to_Cell_rden[34] <= 1'b0;
					reg_FSM_to_Cell_rden[35] <= 1'b0;
					reg_FSM_to_Cell_rden[36] <= 1'b0;
					reg_FSM_to_Cell_rden[37] <= 1'b0;
					reg_FSM_to_Cell_rden[38] <= 1'b0;
					reg_FSM_to_Cell_rden[39] <= 1'b0;
					reg_FSM_to_Cell_rden[40] <= 1'b0;
					reg_FSM_to_Cell_rden[41] <= 1'b0;
					reg_FSM_to_Cell_rden[42] <= 1'b0;
					reg_FSM_to_Cell_rden[43] <= 1'b0;
					reg_FSM_to_Cell_rden[44] <= 1'b0;
					reg_FSM_to_Cell_rden[45] <= 1'b0;
					reg_FSM_to_Cell_rden[46] <= 1'b0;
					reg_FSM_to_Cell_rden[47] <= 1'b0;
					reg_FSM_to_Cell_rden[48] <= 1'b0;
					reg_FSM_to_Cell_rden[49] <= 1'b0;
					reg_FSM_to_Cell_rden[50] <= 1'b0;
					reg_FSM_to_Cell_rden[51] <= 1'b0;
					reg_FSM_to_Cell_rden[52] <= 1'b0;
					reg_FSM_to_Cell_rden[53] <= 1'b0;
					reg_FSM_to_Cell_rden[54] <= 1'b0;
					reg_FSM_to_Cell_rden[55] <= 1'b0;
					reg_FSM_to_Cell_rden[56] <= 1'b0;
					reg_FSM_to_Cell_rden[57] <= 1'b0;
					reg_FSM_to_Cell_rden[58] <= 1'b0;
					reg_FSM_to_Cell_rden[59] <= 1'b0;
					reg_FSM_to_Cell_rden[60] <= 1'b0;
					reg_FSM_to_Cell_rden[61] <= 1'b0;
					reg_FSM_to_Cell_rden[62] <= 1'b0;
					reg_FSM_to_Cell_rden[63] <= 1'b0;
					end
				else
					begin
					reg_FSM_to_Cell_rden[TOTAL_CELL_NUM-1:0] <= 0;
					end
				end
			2:
				begin
				reg_to_force_cache_LJ_Force_Z[1*DATA_WIDTH-1:0*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[2*DATA_WIDTH-1:1*DATA_WIDTH] <= ref_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[3*DATA_WIDTH-1:2*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[4*DATA_WIDTH-1:3*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[5*DATA_WIDTH-1:4*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[6*DATA_WIDTH-1:5*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[7*DATA_WIDTH-1:6*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[8*DATA_WIDTH-1:7*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[9*DATA_WIDTH-1:8*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[10*DATA_WIDTH-1:9*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[11*DATA_WIDTH-1:10*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[12*DATA_WIDTH-1:11*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[13*DATA_WIDTH-1:12*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[14*DATA_WIDTH-1:13*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[15*DATA_WIDTH-1:14*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[16*DATA_WIDTH-1:15*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[17*DATA_WIDTH-1:16*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[18*DATA_WIDTH-1:17*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[19*DATA_WIDTH-1:18*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[20*DATA_WIDTH-1:19*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[21*DATA_WIDTH-1:20*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[22*DATA_WIDTH-1:21*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[23*DATA_WIDTH-1:22*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[24*DATA_WIDTH-1:23*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[25*DATA_WIDTH-1:24*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[26*DATA_WIDTH-1:25*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[27*DATA_WIDTH-1:26*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[28*DATA_WIDTH-1:27*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[29*DATA_WIDTH-1:28*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[30*DATA_WIDTH-1:29*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[31*DATA_WIDTH-1:30*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[32*DATA_WIDTH-1:31*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[33*DATA_WIDTH-1:32*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[34*DATA_WIDTH-1:33*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[35*DATA_WIDTH-1:34*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[36*DATA_WIDTH-1:35*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[37*DATA_WIDTH-1:36*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[38*DATA_WIDTH-1:37*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[39*DATA_WIDTH-1:38*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[40*DATA_WIDTH-1:39*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[41*DATA_WIDTH-1:40*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[42*DATA_WIDTH-1:41*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[43*DATA_WIDTH-1:42*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[44*DATA_WIDTH-1:43*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[45*DATA_WIDTH-1:44*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[46*DATA_WIDTH-1:45*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[47*DATA_WIDTH-1:46*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[48*DATA_WIDTH-1:47*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[49*DATA_WIDTH-1:48*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[50*DATA_WIDTH-1:49*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[51*DATA_WIDTH-1:50*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[52*DATA_WIDTH-1:51*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[53*DATA_WIDTH-1:52*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[54*DATA_WIDTH-1:53*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[55*DATA_WIDTH-1:54*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[56*DATA_WIDTH-1:55*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[57*DATA_WIDTH-1:56*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[58*DATA_WIDTH-1:57*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[59*DATA_WIDTH-1:58*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[60*DATA_WIDTH-1:59*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[61*DATA_WIDTH-1:60*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[62*DATA_WIDTH-1:61*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[63*DATA_WIDTH-1:62*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[64*DATA_WIDTH-1:63*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[1*DATA_WIDTH-1:0*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[2*DATA_WIDTH-1:1*DATA_WIDTH] <= ref_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[3*DATA_WIDTH-1:2*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[4*DATA_WIDTH-1:3*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[5*DATA_WIDTH-1:4*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[6*DATA_WIDTH-1:5*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[7*DATA_WIDTH-1:6*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[8*DATA_WIDTH-1:7*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[9*DATA_WIDTH-1:8*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[10*DATA_WIDTH-1:9*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[11*DATA_WIDTH-1:10*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[12*DATA_WIDTH-1:11*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[13*DATA_WIDTH-1:12*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[14*DATA_WIDTH-1:13*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[15*DATA_WIDTH-1:14*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[16*DATA_WIDTH-1:15*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[17*DATA_WIDTH-1:16*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[18*DATA_WIDTH-1:17*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[19*DATA_WIDTH-1:18*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[20*DATA_WIDTH-1:19*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[21*DATA_WIDTH-1:20*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[22*DATA_WIDTH-1:21*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[23*DATA_WIDTH-1:22*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[24*DATA_WIDTH-1:23*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[25*DATA_WIDTH-1:24*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[26*DATA_WIDTH-1:25*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[27*DATA_WIDTH-1:26*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[28*DATA_WIDTH-1:27*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[29*DATA_WIDTH-1:28*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[30*DATA_WIDTH-1:29*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[31*DATA_WIDTH-1:30*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[32*DATA_WIDTH-1:31*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[33*DATA_WIDTH-1:32*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[34*DATA_WIDTH-1:33*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[35*DATA_WIDTH-1:34*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[36*DATA_WIDTH-1:35*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[37*DATA_WIDTH-1:36*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[38*DATA_WIDTH-1:37*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[39*DATA_WIDTH-1:38*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[40*DATA_WIDTH-1:39*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[41*DATA_WIDTH-1:40*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[42*DATA_WIDTH-1:41*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[43*DATA_WIDTH-1:42*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[44*DATA_WIDTH-1:43*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[45*DATA_WIDTH-1:44*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[46*DATA_WIDTH-1:45*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[47*DATA_WIDTH-1:46*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[48*DATA_WIDTH-1:47*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[49*DATA_WIDTH-1:48*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[50*DATA_WIDTH-1:49*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[51*DATA_WIDTH-1:50*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[52*DATA_WIDTH-1:51*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[53*DATA_WIDTH-1:52*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[54*DATA_WIDTH-1:53*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[55*DATA_WIDTH-1:54*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[56*DATA_WIDTH-1:55*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[57*DATA_WIDTH-1:56*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[58*DATA_WIDTH-1:57*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[59*DATA_WIDTH-1:58*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[60*DATA_WIDTH-1:59*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[61*DATA_WIDTH-1:60*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[62*DATA_WIDTH-1:61*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[63*DATA_WIDTH-1:62*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[64*DATA_WIDTH-1:63*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[1*DATA_WIDTH-1:0*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[2*DATA_WIDTH-1:1*DATA_WIDTH] <= ref_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[3*DATA_WIDTH-1:2*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[4*DATA_WIDTH-1:3*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[5*DATA_WIDTH-1:4*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[6*DATA_WIDTH-1:5*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[7*DATA_WIDTH-1:6*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[8*DATA_WIDTH-1:7*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[9*DATA_WIDTH-1:8*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[10*DATA_WIDTH-1:9*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[11*DATA_WIDTH-1:10*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[12*DATA_WIDTH-1:11*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[13*DATA_WIDTH-1:12*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[14*DATA_WIDTH-1:13*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[15*DATA_WIDTH-1:14*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[16*DATA_WIDTH-1:15*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[17*DATA_WIDTH-1:16*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[18*DATA_WIDTH-1:17*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[19*DATA_WIDTH-1:18*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[20*DATA_WIDTH-1:19*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[21*DATA_WIDTH-1:20*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[22*DATA_WIDTH-1:21*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[23*DATA_WIDTH-1:22*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[24*DATA_WIDTH-1:23*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[25*DATA_WIDTH-1:24*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[26*DATA_WIDTH-1:25*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[27*DATA_WIDTH-1:26*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[28*DATA_WIDTH-1:27*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[29*DATA_WIDTH-1:28*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[30*DATA_WIDTH-1:29*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[31*DATA_WIDTH-1:30*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[32*DATA_WIDTH-1:31*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[33*DATA_WIDTH-1:32*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[34*DATA_WIDTH-1:33*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[35*DATA_WIDTH-1:34*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[36*DATA_WIDTH-1:35*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[37*DATA_WIDTH-1:36*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[38*DATA_WIDTH-1:37*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[39*DATA_WIDTH-1:38*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[40*DATA_WIDTH-1:39*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[41*DATA_WIDTH-1:40*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[42*DATA_WIDTH-1:41*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[43*DATA_WIDTH-1:42*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[44*DATA_WIDTH-1:43*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[45*DATA_WIDTH-1:44*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[46*DATA_WIDTH-1:45*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[47*DATA_WIDTH-1:46*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[48*DATA_WIDTH-1:47*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[49*DATA_WIDTH-1:48*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[50*DATA_WIDTH-1:49*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[51*DATA_WIDTH-1:50*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[52*DATA_WIDTH-1:51*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[53*DATA_WIDTH-1:52*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[54*DATA_WIDTH-1:53*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[55*DATA_WIDTH-1:54*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[56*DATA_WIDTH-1:55*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[57*DATA_WIDTH-1:56*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[58*DATA_WIDTH-1:57*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[59*DATA_WIDTH-1:58*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[60*DATA_WIDTH-1:59*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[61*DATA_WIDTH-1:60*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[62*DATA_WIDTH-1:61*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[63*DATA_WIDTH-1:62*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[64*DATA_WIDTH-1:63*DATA_WIDTH] <= 0;
				reg_to_force_cache_particle_id[1*PARTICLE_ID_WIDTH-1:0*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[2*PARTICLE_ID_WIDTH-1:1*PARTICLE_ID_WIDTH] <= ref_particle_id_1_1;
				reg_to_force_cache_particle_id[3*PARTICLE_ID_WIDTH-1:2*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[4*PARTICLE_ID_WIDTH-1:3*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[5*PARTICLE_ID_WIDTH-1:4*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[6*PARTICLE_ID_WIDTH-1:5*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[7*PARTICLE_ID_WIDTH-1:6*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[8*PARTICLE_ID_WIDTH-1:7*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[9*PARTICLE_ID_WIDTH-1:8*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[10*PARTICLE_ID_WIDTH-1:9*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[11*PARTICLE_ID_WIDTH-1:10*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[12*PARTICLE_ID_WIDTH-1:11*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[13*PARTICLE_ID_WIDTH-1:12*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[14*PARTICLE_ID_WIDTH-1:13*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[15*PARTICLE_ID_WIDTH-1:14*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[16*PARTICLE_ID_WIDTH-1:15*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[17*PARTICLE_ID_WIDTH-1:16*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[18*PARTICLE_ID_WIDTH-1:17*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[19*PARTICLE_ID_WIDTH-1:18*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[20*PARTICLE_ID_WIDTH-1:19*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[21*PARTICLE_ID_WIDTH-1:20*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[22*PARTICLE_ID_WIDTH-1:21*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[23*PARTICLE_ID_WIDTH-1:22*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[24*PARTICLE_ID_WIDTH-1:23*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[25*PARTICLE_ID_WIDTH-1:24*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[26*PARTICLE_ID_WIDTH-1:25*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[27*PARTICLE_ID_WIDTH-1:26*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[28*PARTICLE_ID_WIDTH-1:27*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[29*PARTICLE_ID_WIDTH-1:28*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[30*PARTICLE_ID_WIDTH-1:29*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[31*PARTICLE_ID_WIDTH-1:30*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[32*PARTICLE_ID_WIDTH-1:31*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[33*PARTICLE_ID_WIDTH-1:32*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[34*PARTICLE_ID_WIDTH-1:33*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[35*PARTICLE_ID_WIDTH-1:34*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[36*PARTICLE_ID_WIDTH-1:35*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[37*PARTICLE_ID_WIDTH-1:36*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[38*PARTICLE_ID_WIDTH-1:37*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[39*PARTICLE_ID_WIDTH-1:38*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[40*PARTICLE_ID_WIDTH-1:39*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[41*PARTICLE_ID_WIDTH-1:40*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[42*PARTICLE_ID_WIDTH-1:41*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[43*PARTICLE_ID_WIDTH-1:42*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[44*PARTICLE_ID_WIDTH-1:43*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[45*PARTICLE_ID_WIDTH-1:44*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[46*PARTICLE_ID_WIDTH-1:45*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[47*PARTICLE_ID_WIDTH-1:46*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[48*PARTICLE_ID_WIDTH-1:47*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[49*PARTICLE_ID_WIDTH-1:48*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[50*PARTICLE_ID_WIDTH-1:49*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[51*PARTICLE_ID_WIDTH-1:50*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[52*PARTICLE_ID_WIDTH-1:51*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[53*PARTICLE_ID_WIDTH-1:52*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[54*PARTICLE_ID_WIDTH-1:53*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[55*PARTICLE_ID_WIDTH-1:54*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[56*PARTICLE_ID_WIDTH-1:55*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[57*PARTICLE_ID_WIDTH-1:56*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[58*PARTICLE_ID_WIDTH-1:57*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[59*PARTICLE_ID_WIDTH-1:58*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[60*PARTICLE_ID_WIDTH-1:59*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[61*PARTICLE_ID_WIDTH-1:60*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[62*PARTICLE_ID_WIDTH-1:61*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[63*PARTICLE_ID_WIDTH-1:62*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[64*PARTICLE_ID_WIDTH-1:63*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_partial_force_valid[0] <= 1'b0;
				reg_to_force_cache_partial_force_valid[1] <= ref_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[2] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[3] <= 1'b0;
				reg_to_force_cache_partial_force_valid[4] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[5] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[6] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[7] <= 1'b0;
				reg_to_force_cache_partial_force_valid[8] <= 1'b0;
				reg_to_force_cache_partial_force_valid[9] <= 1'b0;
				reg_to_force_cache_partial_force_valid[10] <= 1'b0;
				reg_to_force_cache_partial_force_valid[11] <= 1'b0;
				reg_to_force_cache_partial_force_valid[12] <= 1'b0;
				reg_to_force_cache_partial_force_valid[13] <= 1'b0;
				reg_to_force_cache_partial_force_valid[14] <= 1'b0;
				reg_to_force_cache_partial_force_valid[15] <= 1'b0;
				reg_to_force_cache_partial_force_valid[16] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[17] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[18] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[19] <= 1'b0;
				reg_to_force_cache_partial_force_valid[20] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[21] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[22] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[23] <= 1'b0;
				reg_to_force_cache_partial_force_valid[24] <= 1'b0;
				reg_to_force_cache_partial_force_valid[25] <= 1'b0;
				reg_to_force_cache_partial_force_valid[26] <= 1'b0;
				reg_to_force_cache_partial_force_valid[27] <= 1'b0;
				reg_to_force_cache_partial_force_valid[28] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[29] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[30] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[31] <= 1'b0;
				reg_to_force_cache_partial_force_valid[32] <= 1'b0;
				reg_to_force_cache_partial_force_valid[33] <= 1'b0;
				reg_to_force_cache_partial_force_valid[34] <= 1'b0;
				reg_to_force_cache_partial_force_valid[35] <= 1'b0;
				reg_to_force_cache_partial_force_valid[36] <= 1'b0;
				reg_to_force_cache_partial_force_valid[37] <= 1'b0;
				reg_to_force_cache_partial_force_valid[38] <= 1'b0;
				reg_to_force_cache_partial_force_valid[39] <= 1'b0;
				reg_to_force_cache_partial_force_valid[40] <= 1'b0;
				reg_to_force_cache_partial_force_valid[41] <= 1'b0;
				reg_to_force_cache_partial_force_valid[42] <= 1'b0;
				reg_to_force_cache_partial_force_valid[43] <= 1'b0;
				reg_to_force_cache_partial_force_valid[44] <= 1'b0;
				reg_to_force_cache_partial_force_valid[45] <= 1'b0;
				reg_to_force_cache_partial_force_valid[46] <= 1'b0;
				reg_to_force_cache_partial_force_valid[47] <= 1'b0;
				reg_to_force_cache_partial_force_valid[48] <= 1'b0;
				reg_to_force_cache_partial_force_valid[49] <= 1'b0;
				reg_to_force_cache_partial_force_valid[50] <= 1'b0;
				reg_to_force_cache_partial_force_valid[51] <= 1'b0;
				reg_to_force_cache_partial_force_valid[52] <= 1'b0;
				reg_to_force_cache_partial_force_valid[53] <= 1'b0;
				reg_to_force_cache_partial_force_valid[54] <= 1'b0;
				reg_to_force_cache_partial_force_valid[55] <= 1'b0;
				reg_to_force_cache_partial_force_valid[56] <= 1'b0;
				reg_to_force_cache_partial_force_valid[57] <= 1'b0;
				reg_to_force_cache_partial_force_valid[58] <= 1'b0;
				reg_to_force_cache_partial_force_valid[59] <= 1'b0;
				reg_to_force_cache_partial_force_valid[60] <= 1'b0;
				reg_to_force_cache_partial_force_valid[61] <= 1'b0;
				reg_to_force_cache_partial_force_valid[62] <= 1'b0;
				reg_to_force_cache_partial_force_valid[63] <= 1'b0;
				reg_cells_to_pipeline_1_1 <= 	{
														Position_Cache_readout_position[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH],
														Position_Cache_readout_position[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH],
														Position_Cache_readout_position[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH],
														Position_Cache_readout_position[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH],
														Position_Cache_readout_position[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH],
														Position_Cache_readout_position[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH],
														Position_Cache_readout_position[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH],
														Position_Cache_readout_position[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH],
														Position_Cache_readout_position[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH],
														Position_Cache_readout_position[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH],
														Position_Cache_readout_position[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH],
														Position_Cache_readout_position[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH],
														Position_Cache_readout_position[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH],
														Position_Cache_readout_position[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH]
														};
				reg_FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[15*CELL_ADDR_WIDTH-1:14*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[16*CELL_ADDR_WIDTH-1:15*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[17*CELL_ADDR_WIDTH-1:16*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[18*CELL_ADDR_WIDTH-1:17*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[19*CELL_ADDR_WIDTH-1:18*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[20*CELL_ADDR_WIDTH-1:19*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[21*CELL_ADDR_WIDTH-1:20*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[22*CELL_ADDR_WIDTH-1:21*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[23*CELL_ADDR_WIDTH-1:22*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[24*CELL_ADDR_WIDTH-1:23*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[25*CELL_ADDR_WIDTH-1:24*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[26*CELL_ADDR_WIDTH-1:25*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[27*CELL_ADDR_WIDTH-1:26*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[28*CELL_ADDR_WIDTH-1:27*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[29*CELL_ADDR_WIDTH-1:28*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[30*CELL_ADDR_WIDTH-1:29*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[31*CELL_ADDR_WIDTH-1:30*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[32*CELL_ADDR_WIDTH-1:31*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[33*CELL_ADDR_WIDTH-1:32*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[34*CELL_ADDR_WIDTH-1:33*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[35*CELL_ADDR_WIDTH-1:34*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[36*CELL_ADDR_WIDTH-1:35*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[37*CELL_ADDR_WIDTH-1:36*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[38*CELL_ADDR_WIDTH-1:37*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[39*CELL_ADDR_WIDTH-1:38*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[40*CELL_ADDR_WIDTH-1:39*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[41*CELL_ADDR_WIDTH-1:40*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[42*CELL_ADDR_WIDTH-1:41*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[43*CELL_ADDR_WIDTH-1:42*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[44*CELL_ADDR_WIDTH-1:43*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[45*CELL_ADDR_WIDTH-1:44*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[46*CELL_ADDR_WIDTH-1:45*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[47*CELL_ADDR_WIDTH-1:46*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[48*CELL_ADDR_WIDTH-1:47*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[49*CELL_ADDR_WIDTH-1:48*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[50*CELL_ADDR_WIDTH-1:49*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[51*CELL_ADDR_WIDTH-1:50*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[52*CELL_ADDR_WIDTH-1:51*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[53*CELL_ADDR_WIDTH-1:52*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[54*CELL_ADDR_WIDTH-1:53*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[55*CELL_ADDR_WIDTH-1:54*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[56*CELL_ADDR_WIDTH-1:55*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[57*CELL_ADDR_WIDTH-1:56*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[58*CELL_ADDR_WIDTH-1:57*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[59*CELL_ADDR_WIDTH-1:58*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[60*CELL_ADDR_WIDTH-1:59*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[61*CELL_ADDR_WIDTH-1:60*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[62*CELL_ADDR_WIDTH-1:61*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[63*CELL_ADDR_WIDTH-1:62*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[64*CELL_ADDR_WIDTH-1:63*CELL_ADDR_WIDTH] <= 0;
				if (FSM_to_Cell_rden_1_1)
					begin
					reg_FSM_to_Cell_rden[0] <= 1'b0;
					reg_FSM_to_Cell_rden[1] <= 1'b1;
					reg_FSM_to_Cell_rden[2] <= 1'b1;
					reg_FSM_to_Cell_rden[3] <= 1'b0;
					reg_FSM_to_Cell_rden[4] <= 1'b1;
					reg_FSM_to_Cell_rden[5] <= 1'b1;
					reg_FSM_to_Cell_rden[6] <= 1'b1;
					reg_FSM_to_Cell_rden[7] <= 1'b0;
					reg_FSM_to_Cell_rden[8] <= 1'b0;
					reg_FSM_to_Cell_rden[9] <= 1'b0;
					reg_FSM_to_Cell_rden[10] <= 1'b0;
					reg_FSM_to_Cell_rden[11] <= 1'b0;
					reg_FSM_to_Cell_rden[12] <= 1'b0;
					reg_FSM_to_Cell_rden[13] <= 1'b0;
					reg_FSM_to_Cell_rden[14] <= 1'b0;
					reg_FSM_to_Cell_rden[15] <= 1'b0;
					reg_FSM_to_Cell_rden[16] <= 1'b1;
					reg_FSM_to_Cell_rden[17] <= 1'b1;
					reg_FSM_to_Cell_rden[18] <= 1'b1;
					reg_FSM_to_Cell_rden[19] <= 1'b0;
					reg_FSM_to_Cell_rden[20] <= 1'b1;
					reg_FSM_to_Cell_rden[21] <= 1'b1;
					reg_FSM_to_Cell_rden[22] <= 1'b1;
					reg_FSM_to_Cell_rden[23] <= 1'b0;
					reg_FSM_to_Cell_rden[24] <= 1'b0;
					reg_FSM_to_Cell_rden[25] <= 1'b0;
					reg_FSM_to_Cell_rden[26] <= 1'b0;
					reg_FSM_to_Cell_rden[27] <= 1'b0;
					reg_FSM_to_Cell_rden[28] <= 1'b1;
					reg_FSM_to_Cell_rden[29] <= 1'b1;
					reg_FSM_to_Cell_rden[30] <= 1'b1;
					reg_FSM_to_Cell_rden[31] <= 1'b0;
					reg_FSM_to_Cell_rden[32] <= 1'b0;
					reg_FSM_to_Cell_rden[33] <= 1'b0;
					reg_FSM_to_Cell_rden[34] <= 1'b0;
					reg_FSM_to_Cell_rden[35] <= 1'b0;
					reg_FSM_to_Cell_rden[36] <= 1'b0;
					reg_FSM_to_Cell_rden[37] <= 1'b0;
					reg_FSM_to_Cell_rden[38] <= 1'b0;
					reg_FSM_to_Cell_rden[39] <= 1'b0;
					reg_FSM_to_Cell_rden[40] <= 1'b0;
					reg_FSM_to_Cell_rden[41] <= 1'b0;
					reg_FSM_to_Cell_rden[42] <= 1'b0;
					reg_FSM_to_Cell_rden[43] <= 1'b0;
					reg_FSM_to_Cell_rden[44] <= 1'b0;
					reg_FSM_to_Cell_rden[45] <= 1'b0;
					reg_FSM_to_Cell_rden[46] <= 1'b0;
					reg_FSM_to_Cell_rden[47] <= 1'b0;
					reg_FSM_to_Cell_rden[48] <= 1'b0;
					reg_FSM_to_Cell_rden[49] <= 1'b0;
					reg_FSM_to_Cell_rden[50] <= 1'b0;
					reg_FSM_to_Cell_rden[51] <= 1'b0;
					reg_FSM_to_Cell_rden[52] <= 1'b0;
					reg_FSM_to_Cell_rden[53] <= 1'b0;
					reg_FSM_to_Cell_rden[54] <= 1'b0;
					reg_FSM_to_Cell_rden[55] <= 1'b0;
					reg_FSM_to_Cell_rden[56] <= 1'b0;
					reg_FSM_to_Cell_rden[57] <= 1'b0;
					reg_FSM_to_Cell_rden[58] <= 1'b0;
					reg_FSM_to_Cell_rden[59] <= 1'b0;
					reg_FSM_to_Cell_rden[60] <= 1'b0;
					reg_FSM_to_Cell_rden[61] <= 1'b0;
					reg_FSM_to_Cell_rden[62] <= 1'b0;
					reg_FSM_to_Cell_rden[63] <= 1'b0;
					end
				else
					begin
					reg_FSM_to_Cell_rden[TOTAL_CELL_NUM-1:0] <= 0;
					end
				end
			3:
				begin
				reg_to_force_cache_LJ_Force_Z[1*DATA_WIDTH-1:0*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[2*DATA_WIDTH-1:1*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[3*DATA_WIDTH-1:2*DATA_WIDTH] <= ref_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[4*DATA_WIDTH-1:3*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[5*DATA_WIDTH-1:4*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[6*DATA_WIDTH-1:5*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[7*DATA_WIDTH-1:6*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[8*DATA_WIDTH-1:7*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[9*DATA_WIDTH-1:8*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[10*DATA_WIDTH-1:9*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[11*DATA_WIDTH-1:10*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[12*DATA_WIDTH-1:11*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[13*DATA_WIDTH-1:12*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[14*DATA_WIDTH-1:13*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[15*DATA_WIDTH-1:14*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[16*DATA_WIDTH-1:15*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[17*DATA_WIDTH-1:16*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[18*DATA_WIDTH-1:17*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[19*DATA_WIDTH-1:18*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[20*DATA_WIDTH-1:19*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[21*DATA_WIDTH-1:20*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[22*DATA_WIDTH-1:21*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[23*DATA_WIDTH-1:22*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[24*DATA_WIDTH-1:23*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[25*DATA_WIDTH-1:24*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[26*DATA_WIDTH-1:25*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[27*DATA_WIDTH-1:26*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[28*DATA_WIDTH-1:27*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[29*DATA_WIDTH-1:28*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[30*DATA_WIDTH-1:29*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[31*DATA_WIDTH-1:30*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[32*DATA_WIDTH-1:31*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[33*DATA_WIDTH-1:32*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[34*DATA_WIDTH-1:33*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[35*DATA_WIDTH-1:34*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[36*DATA_WIDTH-1:35*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[37*DATA_WIDTH-1:36*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[38*DATA_WIDTH-1:37*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[39*DATA_WIDTH-1:38*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[40*DATA_WIDTH-1:39*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[41*DATA_WIDTH-1:40*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[42*DATA_WIDTH-1:41*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[43*DATA_WIDTH-1:42*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[44*DATA_WIDTH-1:43*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[45*DATA_WIDTH-1:44*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[46*DATA_WIDTH-1:45*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[47*DATA_WIDTH-1:46*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[48*DATA_WIDTH-1:47*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[49*DATA_WIDTH-1:48*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[50*DATA_WIDTH-1:49*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[51*DATA_WIDTH-1:50*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[52*DATA_WIDTH-1:51*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[53*DATA_WIDTH-1:52*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[54*DATA_WIDTH-1:53*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[55*DATA_WIDTH-1:54*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[56*DATA_WIDTH-1:55*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[57*DATA_WIDTH-1:56*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[58*DATA_WIDTH-1:57*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[59*DATA_WIDTH-1:58*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[60*DATA_WIDTH-1:59*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[61*DATA_WIDTH-1:60*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[62*DATA_WIDTH-1:61*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[63*DATA_WIDTH-1:62*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[64*DATA_WIDTH-1:63*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[1*DATA_WIDTH-1:0*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[2*DATA_WIDTH-1:1*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[3*DATA_WIDTH-1:2*DATA_WIDTH] <= ref_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[4*DATA_WIDTH-1:3*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[5*DATA_WIDTH-1:4*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[6*DATA_WIDTH-1:5*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[7*DATA_WIDTH-1:6*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[8*DATA_WIDTH-1:7*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[9*DATA_WIDTH-1:8*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[10*DATA_WIDTH-1:9*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[11*DATA_WIDTH-1:10*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[12*DATA_WIDTH-1:11*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[13*DATA_WIDTH-1:12*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[14*DATA_WIDTH-1:13*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[15*DATA_WIDTH-1:14*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[16*DATA_WIDTH-1:15*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[17*DATA_WIDTH-1:16*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[18*DATA_WIDTH-1:17*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[19*DATA_WIDTH-1:18*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[20*DATA_WIDTH-1:19*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[21*DATA_WIDTH-1:20*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[22*DATA_WIDTH-1:21*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[23*DATA_WIDTH-1:22*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[24*DATA_WIDTH-1:23*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[25*DATA_WIDTH-1:24*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[26*DATA_WIDTH-1:25*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[27*DATA_WIDTH-1:26*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[28*DATA_WIDTH-1:27*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[29*DATA_WIDTH-1:28*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[30*DATA_WIDTH-1:29*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[31*DATA_WIDTH-1:30*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[32*DATA_WIDTH-1:31*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[33*DATA_WIDTH-1:32*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[34*DATA_WIDTH-1:33*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[35*DATA_WIDTH-1:34*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[36*DATA_WIDTH-1:35*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[37*DATA_WIDTH-1:36*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[38*DATA_WIDTH-1:37*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[39*DATA_WIDTH-1:38*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[40*DATA_WIDTH-1:39*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[41*DATA_WIDTH-1:40*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[42*DATA_WIDTH-1:41*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[43*DATA_WIDTH-1:42*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[44*DATA_WIDTH-1:43*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[45*DATA_WIDTH-1:44*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[46*DATA_WIDTH-1:45*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[47*DATA_WIDTH-1:46*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[48*DATA_WIDTH-1:47*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[49*DATA_WIDTH-1:48*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[50*DATA_WIDTH-1:49*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[51*DATA_WIDTH-1:50*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[52*DATA_WIDTH-1:51*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[53*DATA_WIDTH-1:52*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[54*DATA_WIDTH-1:53*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[55*DATA_WIDTH-1:54*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[56*DATA_WIDTH-1:55*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[57*DATA_WIDTH-1:56*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[58*DATA_WIDTH-1:57*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[59*DATA_WIDTH-1:58*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[60*DATA_WIDTH-1:59*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[61*DATA_WIDTH-1:60*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[62*DATA_WIDTH-1:61*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[63*DATA_WIDTH-1:62*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[64*DATA_WIDTH-1:63*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[1*DATA_WIDTH-1:0*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[2*DATA_WIDTH-1:1*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[3*DATA_WIDTH-1:2*DATA_WIDTH] <= ref_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[4*DATA_WIDTH-1:3*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[5*DATA_WIDTH-1:4*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[6*DATA_WIDTH-1:5*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[7*DATA_WIDTH-1:6*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[8*DATA_WIDTH-1:7*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[9*DATA_WIDTH-1:8*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[10*DATA_WIDTH-1:9*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[11*DATA_WIDTH-1:10*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[12*DATA_WIDTH-1:11*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[13*DATA_WIDTH-1:12*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[14*DATA_WIDTH-1:13*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[15*DATA_WIDTH-1:14*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[16*DATA_WIDTH-1:15*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[17*DATA_WIDTH-1:16*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[18*DATA_WIDTH-1:17*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[19*DATA_WIDTH-1:18*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[20*DATA_WIDTH-1:19*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[21*DATA_WIDTH-1:20*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[22*DATA_WIDTH-1:21*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[23*DATA_WIDTH-1:22*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[24*DATA_WIDTH-1:23*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[25*DATA_WIDTH-1:24*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[26*DATA_WIDTH-1:25*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[27*DATA_WIDTH-1:26*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[28*DATA_WIDTH-1:27*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[29*DATA_WIDTH-1:28*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[30*DATA_WIDTH-1:29*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[31*DATA_WIDTH-1:30*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[32*DATA_WIDTH-1:31*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[33*DATA_WIDTH-1:32*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[34*DATA_WIDTH-1:33*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[35*DATA_WIDTH-1:34*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[36*DATA_WIDTH-1:35*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[37*DATA_WIDTH-1:36*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[38*DATA_WIDTH-1:37*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[39*DATA_WIDTH-1:38*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[40*DATA_WIDTH-1:39*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[41*DATA_WIDTH-1:40*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[42*DATA_WIDTH-1:41*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[43*DATA_WIDTH-1:42*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[44*DATA_WIDTH-1:43*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[45*DATA_WIDTH-1:44*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[46*DATA_WIDTH-1:45*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[47*DATA_WIDTH-1:46*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[48*DATA_WIDTH-1:47*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[49*DATA_WIDTH-1:48*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[50*DATA_WIDTH-1:49*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[51*DATA_WIDTH-1:50*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[52*DATA_WIDTH-1:51*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[53*DATA_WIDTH-1:52*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[54*DATA_WIDTH-1:53*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[55*DATA_WIDTH-1:54*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[56*DATA_WIDTH-1:55*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[57*DATA_WIDTH-1:56*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[58*DATA_WIDTH-1:57*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[59*DATA_WIDTH-1:58*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[60*DATA_WIDTH-1:59*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[61*DATA_WIDTH-1:60*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[62*DATA_WIDTH-1:61*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[63*DATA_WIDTH-1:62*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[64*DATA_WIDTH-1:63*DATA_WIDTH] <= 0;
				reg_to_force_cache_particle_id[1*PARTICLE_ID_WIDTH-1:0*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[2*PARTICLE_ID_WIDTH-1:1*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[3*PARTICLE_ID_WIDTH-1:2*PARTICLE_ID_WIDTH] <= ref_particle_id_1_1;
				reg_to_force_cache_particle_id[4*PARTICLE_ID_WIDTH-1:3*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[5*PARTICLE_ID_WIDTH-1:4*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[6*PARTICLE_ID_WIDTH-1:5*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[7*PARTICLE_ID_WIDTH-1:6*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[8*PARTICLE_ID_WIDTH-1:7*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[9*PARTICLE_ID_WIDTH-1:8*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[10*PARTICLE_ID_WIDTH-1:9*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[11*PARTICLE_ID_WIDTH-1:10*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[12*PARTICLE_ID_WIDTH-1:11*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[13*PARTICLE_ID_WIDTH-1:12*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[14*PARTICLE_ID_WIDTH-1:13*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[15*PARTICLE_ID_WIDTH-1:14*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[16*PARTICLE_ID_WIDTH-1:15*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[17*PARTICLE_ID_WIDTH-1:16*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[18*PARTICLE_ID_WIDTH-1:17*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[19*PARTICLE_ID_WIDTH-1:18*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[20*PARTICLE_ID_WIDTH-1:19*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[21*PARTICLE_ID_WIDTH-1:20*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[22*PARTICLE_ID_WIDTH-1:21*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[23*PARTICLE_ID_WIDTH-1:22*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[24*PARTICLE_ID_WIDTH-1:23*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[25*PARTICLE_ID_WIDTH-1:24*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[26*PARTICLE_ID_WIDTH-1:25*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[27*PARTICLE_ID_WIDTH-1:26*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[28*PARTICLE_ID_WIDTH-1:27*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[29*PARTICLE_ID_WIDTH-1:28*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[30*PARTICLE_ID_WIDTH-1:29*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[31*PARTICLE_ID_WIDTH-1:30*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[32*PARTICLE_ID_WIDTH-1:31*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[33*PARTICLE_ID_WIDTH-1:32*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[34*PARTICLE_ID_WIDTH-1:33*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[35*PARTICLE_ID_WIDTH-1:34*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[36*PARTICLE_ID_WIDTH-1:35*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[37*PARTICLE_ID_WIDTH-1:36*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[38*PARTICLE_ID_WIDTH-1:37*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[39*PARTICLE_ID_WIDTH-1:38*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[40*PARTICLE_ID_WIDTH-1:39*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[41*PARTICLE_ID_WIDTH-1:40*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[42*PARTICLE_ID_WIDTH-1:41*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[43*PARTICLE_ID_WIDTH-1:42*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[44*PARTICLE_ID_WIDTH-1:43*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[45*PARTICLE_ID_WIDTH-1:44*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[46*PARTICLE_ID_WIDTH-1:45*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[47*PARTICLE_ID_WIDTH-1:46*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[48*PARTICLE_ID_WIDTH-1:47*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[49*PARTICLE_ID_WIDTH-1:48*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[50*PARTICLE_ID_WIDTH-1:49*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[51*PARTICLE_ID_WIDTH-1:50*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[52*PARTICLE_ID_WIDTH-1:51*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[53*PARTICLE_ID_WIDTH-1:52*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[54*PARTICLE_ID_WIDTH-1:53*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[55*PARTICLE_ID_WIDTH-1:54*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[56*PARTICLE_ID_WIDTH-1:55*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[57*PARTICLE_ID_WIDTH-1:56*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[58*PARTICLE_ID_WIDTH-1:57*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[59*PARTICLE_ID_WIDTH-1:58*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[60*PARTICLE_ID_WIDTH-1:59*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[61*PARTICLE_ID_WIDTH-1:60*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[62*PARTICLE_ID_WIDTH-1:61*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[63*PARTICLE_ID_WIDTH-1:62*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[64*PARTICLE_ID_WIDTH-1:63*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_partial_force_valid[0] <= 1'b0;
				reg_to_force_cache_partial_force_valid[1] <= 1'b0;
				reg_to_force_cache_partial_force_valid[2] <= ref_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[3] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[4] <= 1'b0;
				reg_to_force_cache_partial_force_valid[5] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[6] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[7] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[8] <= 1'b0;
				reg_to_force_cache_partial_force_valid[9] <= 1'b0;
				reg_to_force_cache_partial_force_valid[10] <= 1'b0;
				reg_to_force_cache_partial_force_valid[11] <= 1'b0;
				reg_to_force_cache_partial_force_valid[12] <= 1'b0;
				reg_to_force_cache_partial_force_valid[13] <= 1'b0;
				reg_to_force_cache_partial_force_valid[14] <= 1'b0;
				reg_to_force_cache_partial_force_valid[15] <= 1'b0;
				reg_to_force_cache_partial_force_valid[16] <= 1'b0;
				reg_to_force_cache_partial_force_valid[17] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[18] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[19] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[20] <= 1'b0;
				reg_to_force_cache_partial_force_valid[21] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[22] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[23] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[24] <= 1'b0;
				reg_to_force_cache_partial_force_valid[25] <= 1'b0;
				reg_to_force_cache_partial_force_valid[26] <= 1'b0;
				reg_to_force_cache_partial_force_valid[27] <= 1'b0;
				reg_to_force_cache_partial_force_valid[28] <= 1'b0;
				reg_to_force_cache_partial_force_valid[29] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[30] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[31] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[32] <= 1'b0;
				reg_to_force_cache_partial_force_valid[33] <= 1'b0;
				reg_to_force_cache_partial_force_valid[34] <= 1'b0;
				reg_to_force_cache_partial_force_valid[35] <= 1'b0;
				reg_to_force_cache_partial_force_valid[36] <= 1'b0;
				reg_to_force_cache_partial_force_valid[37] <= 1'b0;
				reg_to_force_cache_partial_force_valid[38] <= 1'b0;
				reg_to_force_cache_partial_force_valid[39] <= 1'b0;
				reg_to_force_cache_partial_force_valid[40] <= 1'b0;
				reg_to_force_cache_partial_force_valid[41] <= 1'b0;
				reg_to_force_cache_partial_force_valid[42] <= 1'b0;
				reg_to_force_cache_partial_force_valid[43] <= 1'b0;
				reg_to_force_cache_partial_force_valid[44] <= 1'b0;
				reg_to_force_cache_partial_force_valid[45] <= 1'b0;
				reg_to_force_cache_partial_force_valid[46] <= 1'b0;
				reg_to_force_cache_partial_force_valid[47] <= 1'b0;
				reg_to_force_cache_partial_force_valid[48] <= 1'b0;
				reg_to_force_cache_partial_force_valid[49] <= 1'b0;
				reg_to_force_cache_partial_force_valid[50] <= 1'b0;
				reg_to_force_cache_partial_force_valid[51] <= 1'b0;
				reg_to_force_cache_partial_force_valid[52] <= 1'b0;
				reg_to_force_cache_partial_force_valid[53] <= 1'b0;
				reg_to_force_cache_partial_force_valid[54] <= 1'b0;
				reg_to_force_cache_partial_force_valid[55] <= 1'b0;
				reg_to_force_cache_partial_force_valid[56] <= 1'b0;
				reg_to_force_cache_partial_force_valid[57] <= 1'b0;
				reg_to_force_cache_partial_force_valid[58] <= 1'b0;
				reg_to_force_cache_partial_force_valid[59] <= 1'b0;
				reg_to_force_cache_partial_force_valid[60] <= 1'b0;
				reg_to_force_cache_partial_force_valid[61] <= 1'b0;
				reg_to_force_cache_partial_force_valid[62] <= 1'b0;
				reg_to_force_cache_partial_force_valid[63] <= 1'b0;
				reg_cells_to_pipeline_1_1 <= 	{
														Position_Cache_readout_position[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH],
														Position_Cache_readout_position[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH],
														Position_Cache_readout_position[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH],
														Position_Cache_readout_position[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH],
														Position_Cache_readout_position[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH],
														Position_Cache_readout_position[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH],
														Position_Cache_readout_position[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH],
														Position_Cache_readout_position[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH],
														Position_Cache_readout_position[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH],
														Position_Cache_readout_position[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH],
														Position_Cache_readout_position[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH],
														Position_Cache_readout_position[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH],
														Position_Cache_readout_position[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH],
														Position_Cache_readout_position[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH]
														};
				reg_FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[15*CELL_ADDR_WIDTH-1:14*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[16*CELL_ADDR_WIDTH-1:15*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[17*CELL_ADDR_WIDTH-1:16*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[18*CELL_ADDR_WIDTH-1:17*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[19*CELL_ADDR_WIDTH-1:18*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[20*CELL_ADDR_WIDTH-1:19*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[21*CELL_ADDR_WIDTH-1:20*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[22*CELL_ADDR_WIDTH-1:21*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[23*CELL_ADDR_WIDTH-1:22*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[24*CELL_ADDR_WIDTH-1:23*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[25*CELL_ADDR_WIDTH-1:24*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[26*CELL_ADDR_WIDTH-1:25*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[27*CELL_ADDR_WIDTH-1:26*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[28*CELL_ADDR_WIDTH-1:27*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[29*CELL_ADDR_WIDTH-1:28*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[30*CELL_ADDR_WIDTH-1:29*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[31*CELL_ADDR_WIDTH-1:30*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[32*CELL_ADDR_WIDTH-1:31*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[33*CELL_ADDR_WIDTH-1:32*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[34*CELL_ADDR_WIDTH-1:33*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[35*CELL_ADDR_WIDTH-1:34*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[36*CELL_ADDR_WIDTH-1:35*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[37*CELL_ADDR_WIDTH-1:36*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[38*CELL_ADDR_WIDTH-1:37*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[39*CELL_ADDR_WIDTH-1:38*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[40*CELL_ADDR_WIDTH-1:39*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[41*CELL_ADDR_WIDTH-1:40*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[42*CELL_ADDR_WIDTH-1:41*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[43*CELL_ADDR_WIDTH-1:42*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[44*CELL_ADDR_WIDTH-1:43*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[45*CELL_ADDR_WIDTH-1:44*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[46*CELL_ADDR_WIDTH-1:45*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[47*CELL_ADDR_WIDTH-1:46*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[48*CELL_ADDR_WIDTH-1:47*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[49*CELL_ADDR_WIDTH-1:48*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[50*CELL_ADDR_WIDTH-1:49*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[51*CELL_ADDR_WIDTH-1:50*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[52*CELL_ADDR_WIDTH-1:51*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[53*CELL_ADDR_WIDTH-1:52*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[54*CELL_ADDR_WIDTH-1:53*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[55*CELL_ADDR_WIDTH-1:54*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[56*CELL_ADDR_WIDTH-1:55*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[57*CELL_ADDR_WIDTH-1:56*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[58*CELL_ADDR_WIDTH-1:57*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[59*CELL_ADDR_WIDTH-1:58*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[60*CELL_ADDR_WIDTH-1:59*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[61*CELL_ADDR_WIDTH-1:60*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[62*CELL_ADDR_WIDTH-1:61*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[63*CELL_ADDR_WIDTH-1:62*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[64*CELL_ADDR_WIDTH-1:63*CELL_ADDR_WIDTH] <= 0;
				if (FSM_to_Cell_rden_1_1)
					begin
					reg_FSM_to_Cell_rden[0] <= 1'b0;
					reg_FSM_to_Cell_rden[1] <= 1'b0;
					reg_FSM_to_Cell_rden[2] <= 1'b1;
					reg_FSM_to_Cell_rden[3] <= 1'b1;
					reg_FSM_to_Cell_rden[4] <= 1'b0;
					reg_FSM_to_Cell_rden[5] <= 1'b1;
					reg_FSM_to_Cell_rden[6] <= 1'b1;
					reg_FSM_to_Cell_rden[7] <= 1'b1;
					reg_FSM_to_Cell_rden[8] <= 1'b0;
					reg_FSM_to_Cell_rden[9] <= 1'b0;
					reg_FSM_to_Cell_rden[10] <= 1'b0;
					reg_FSM_to_Cell_rden[11] <= 1'b0;
					reg_FSM_to_Cell_rden[12] <= 1'b0;
					reg_FSM_to_Cell_rden[13] <= 1'b0;
					reg_FSM_to_Cell_rden[14] <= 1'b0;
					reg_FSM_to_Cell_rden[15] <= 1'b0;
					reg_FSM_to_Cell_rden[16] <= 1'b0;
					reg_FSM_to_Cell_rden[17] <= 1'b1;
					reg_FSM_to_Cell_rden[18] <= 1'b1;
					reg_FSM_to_Cell_rden[19] <= 1'b1;
					reg_FSM_to_Cell_rden[20] <= 1'b0;
					reg_FSM_to_Cell_rden[21] <= 1'b1;
					reg_FSM_to_Cell_rden[22] <= 1'b1;
					reg_FSM_to_Cell_rden[23] <= 1'b1;
					reg_FSM_to_Cell_rden[24] <= 1'b0;
					reg_FSM_to_Cell_rden[25] <= 1'b0;
					reg_FSM_to_Cell_rden[26] <= 1'b0;
					reg_FSM_to_Cell_rden[27] <= 1'b0;
					reg_FSM_to_Cell_rden[28] <= 1'b0;
					reg_FSM_to_Cell_rden[29] <= 1'b1;
					reg_FSM_to_Cell_rden[30] <= 1'b1;
					reg_FSM_to_Cell_rden[31] <= 1'b1;
					reg_FSM_to_Cell_rden[32] <= 1'b0;
					reg_FSM_to_Cell_rden[33] <= 1'b0;
					reg_FSM_to_Cell_rden[34] <= 1'b0;
					reg_FSM_to_Cell_rden[35] <= 1'b0;
					reg_FSM_to_Cell_rden[36] <= 1'b0;
					reg_FSM_to_Cell_rden[37] <= 1'b0;
					reg_FSM_to_Cell_rden[38] <= 1'b0;
					reg_FSM_to_Cell_rden[39] <= 1'b0;
					reg_FSM_to_Cell_rden[40] <= 1'b0;
					reg_FSM_to_Cell_rden[41] <= 1'b0;
					reg_FSM_to_Cell_rden[42] <= 1'b0;
					reg_FSM_to_Cell_rden[43] <= 1'b0;
					reg_FSM_to_Cell_rden[44] <= 1'b0;
					reg_FSM_to_Cell_rden[45] <= 1'b0;
					reg_FSM_to_Cell_rden[46] <= 1'b0;
					reg_FSM_to_Cell_rden[47] <= 1'b0;
					reg_FSM_to_Cell_rden[48] <= 1'b0;
					reg_FSM_to_Cell_rden[49] <= 1'b0;
					reg_FSM_to_Cell_rden[50] <= 1'b0;
					reg_FSM_to_Cell_rden[51] <= 1'b0;
					reg_FSM_to_Cell_rden[52] <= 1'b0;
					reg_FSM_to_Cell_rden[53] <= 1'b0;
					reg_FSM_to_Cell_rden[54] <= 1'b0;
					reg_FSM_to_Cell_rden[55] <= 1'b0;
					reg_FSM_to_Cell_rden[56] <= 1'b0;
					reg_FSM_to_Cell_rden[57] <= 1'b0;
					reg_FSM_to_Cell_rden[58] <= 1'b0;
					reg_FSM_to_Cell_rden[59] <= 1'b0;
					reg_FSM_to_Cell_rden[60] <= 1'b0;
					reg_FSM_to_Cell_rden[61] <= 1'b0;
					reg_FSM_to_Cell_rden[62] <= 1'b0;
					reg_FSM_to_Cell_rden[63] <= 1'b0;
					end
				else
					begin
					reg_FSM_to_Cell_rden[TOTAL_CELL_NUM-1:0] <= 0;
					end
				end
			4:
				begin
				reg_to_force_cache_LJ_Force_Z[1*DATA_WIDTH-1:0*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[2*DATA_WIDTH-1:1*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[3*DATA_WIDTH-1:2*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[4*DATA_WIDTH-1:3*DATA_WIDTH] <= ref_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[5*DATA_WIDTH-1:4*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[6*DATA_WIDTH-1:5*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[7*DATA_WIDTH-1:6*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[8*DATA_WIDTH-1:7*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[9*DATA_WIDTH-1:8*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[10*DATA_WIDTH-1:9*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[11*DATA_WIDTH-1:10*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[12*DATA_WIDTH-1:11*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[13*DATA_WIDTH-1:12*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[14*DATA_WIDTH-1:13*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[15*DATA_WIDTH-1:14*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[16*DATA_WIDTH-1:15*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[17*DATA_WIDTH-1:16*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[18*DATA_WIDTH-1:17*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[19*DATA_WIDTH-1:18*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[20*DATA_WIDTH-1:19*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[21*DATA_WIDTH-1:20*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[22*DATA_WIDTH-1:21*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[23*DATA_WIDTH-1:22*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[24*DATA_WIDTH-1:23*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[25*DATA_WIDTH-1:24*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[26*DATA_WIDTH-1:25*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[27*DATA_WIDTH-1:26*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[28*DATA_WIDTH-1:27*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[29*DATA_WIDTH-1:28*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[30*DATA_WIDTH-1:29*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[31*DATA_WIDTH-1:30*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[32*DATA_WIDTH-1:31*DATA_WIDTH] <= neighbor_LJ_Force_Z_1_1;
				reg_to_force_cache_LJ_Force_Z[33*DATA_WIDTH-1:32*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[34*DATA_WIDTH-1:33*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[35*DATA_WIDTH-1:34*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[36*DATA_WIDTH-1:35*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[37*DATA_WIDTH-1:36*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[38*DATA_WIDTH-1:37*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[39*DATA_WIDTH-1:38*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[40*DATA_WIDTH-1:39*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[41*DATA_WIDTH-1:40*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[42*DATA_WIDTH-1:41*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[43*DATA_WIDTH-1:42*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[44*DATA_WIDTH-1:43*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[45*DATA_WIDTH-1:44*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[46*DATA_WIDTH-1:45*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[47*DATA_WIDTH-1:46*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[48*DATA_WIDTH-1:47*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[49*DATA_WIDTH-1:48*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[50*DATA_WIDTH-1:49*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[51*DATA_WIDTH-1:50*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[52*DATA_WIDTH-1:51*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[53*DATA_WIDTH-1:52*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[54*DATA_WIDTH-1:53*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[55*DATA_WIDTH-1:54*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[56*DATA_WIDTH-1:55*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[57*DATA_WIDTH-1:56*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[58*DATA_WIDTH-1:57*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[59*DATA_WIDTH-1:58*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[60*DATA_WIDTH-1:59*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[61*DATA_WIDTH-1:60*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[62*DATA_WIDTH-1:61*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[63*DATA_WIDTH-1:62*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Z[64*DATA_WIDTH-1:63*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[1*DATA_WIDTH-1:0*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[2*DATA_WIDTH-1:1*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[3*DATA_WIDTH-1:2*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[4*DATA_WIDTH-1:3*DATA_WIDTH] <= ref_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[5*DATA_WIDTH-1:4*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[6*DATA_WIDTH-1:5*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[7*DATA_WIDTH-1:6*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[8*DATA_WIDTH-1:7*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[9*DATA_WIDTH-1:8*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[10*DATA_WIDTH-1:9*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[11*DATA_WIDTH-1:10*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[12*DATA_WIDTH-1:11*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[13*DATA_WIDTH-1:12*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[14*DATA_WIDTH-1:13*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[15*DATA_WIDTH-1:14*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[16*DATA_WIDTH-1:15*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[17*DATA_WIDTH-1:16*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[18*DATA_WIDTH-1:17*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[19*DATA_WIDTH-1:18*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[20*DATA_WIDTH-1:19*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[21*DATA_WIDTH-1:20*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[22*DATA_WIDTH-1:21*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[23*DATA_WIDTH-1:22*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[24*DATA_WIDTH-1:23*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[25*DATA_WIDTH-1:24*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[26*DATA_WIDTH-1:25*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[27*DATA_WIDTH-1:26*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[28*DATA_WIDTH-1:27*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[29*DATA_WIDTH-1:28*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[30*DATA_WIDTH-1:29*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[31*DATA_WIDTH-1:30*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[32*DATA_WIDTH-1:31*DATA_WIDTH] <= neighbor_LJ_Force_Y_1_1;
				reg_to_force_cache_LJ_Force_Y[33*DATA_WIDTH-1:32*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[34*DATA_WIDTH-1:33*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[35*DATA_WIDTH-1:34*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[36*DATA_WIDTH-1:35*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[37*DATA_WIDTH-1:36*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[38*DATA_WIDTH-1:37*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[39*DATA_WIDTH-1:38*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[40*DATA_WIDTH-1:39*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[41*DATA_WIDTH-1:40*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[42*DATA_WIDTH-1:41*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[43*DATA_WIDTH-1:42*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[44*DATA_WIDTH-1:43*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[45*DATA_WIDTH-1:44*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[46*DATA_WIDTH-1:45*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[47*DATA_WIDTH-1:46*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[48*DATA_WIDTH-1:47*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[49*DATA_WIDTH-1:48*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[50*DATA_WIDTH-1:49*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[51*DATA_WIDTH-1:50*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[52*DATA_WIDTH-1:51*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[53*DATA_WIDTH-1:52*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[54*DATA_WIDTH-1:53*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[55*DATA_WIDTH-1:54*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[56*DATA_WIDTH-1:55*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[57*DATA_WIDTH-1:56*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[58*DATA_WIDTH-1:57*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[59*DATA_WIDTH-1:58*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[60*DATA_WIDTH-1:59*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[61*DATA_WIDTH-1:60*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[62*DATA_WIDTH-1:61*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[63*DATA_WIDTH-1:62*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_Y[64*DATA_WIDTH-1:63*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[1*DATA_WIDTH-1:0*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[2*DATA_WIDTH-1:1*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[3*DATA_WIDTH-1:2*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[4*DATA_WIDTH-1:3*DATA_WIDTH] <= ref_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[5*DATA_WIDTH-1:4*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[6*DATA_WIDTH-1:5*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[7*DATA_WIDTH-1:6*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[8*DATA_WIDTH-1:7*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[9*DATA_WIDTH-1:8*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[10*DATA_WIDTH-1:9*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[11*DATA_WIDTH-1:10*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[12*DATA_WIDTH-1:11*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[13*DATA_WIDTH-1:12*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[14*DATA_WIDTH-1:13*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[15*DATA_WIDTH-1:14*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[16*DATA_WIDTH-1:15*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[17*DATA_WIDTH-1:16*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[18*DATA_WIDTH-1:17*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[19*DATA_WIDTH-1:18*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[20*DATA_WIDTH-1:19*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[21*DATA_WIDTH-1:20*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[22*DATA_WIDTH-1:21*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[23*DATA_WIDTH-1:22*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[24*DATA_WIDTH-1:23*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[25*DATA_WIDTH-1:24*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[26*DATA_WIDTH-1:25*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[27*DATA_WIDTH-1:26*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[28*DATA_WIDTH-1:27*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[29*DATA_WIDTH-1:28*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[30*DATA_WIDTH-1:29*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[31*DATA_WIDTH-1:30*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[32*DATA_WIDTH-1:31*DATA_WIDTH] <= neighbor_LJ_Force_X_1_1;
				reg_to_force_cache_LJ_Force_X[33*DATA_WIDTH-1:32*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[34*DATA_WIDTH-1:33*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[35*DATA_WIDTH-1:34*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[36*DATA_WIDTH-1:35*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[37*DATA_WIDTH-1:36*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[38*DATA_WIDTH-1:37*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[39*DATA_WIDTH-1:38*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[40*DATA_WIDTH-1:39*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[41*DATA_WIDTH-1:40*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[42*DATA_WIDTH-1:41*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[43*DATA_WIDTH-1:42*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[44*DATA_WIDTH-1:43*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[45*DATA_WIDTH-1:44*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[46*DATA_WIDTH-1:45*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[47*DATA_WIDTH-1:46*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[48*DATA_WIDTH-1:47*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[49*DATA_WIDTH-1:48*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[50*DATA_WIDTH-1:49*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[51*DATA_WIDTH-1:50*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[52*DATA_WIDTH-1:51*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[53*DATA_WIDTH-1:52*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[54*DATA_WIDTH-1:53*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[55*DATA_WIDTH-1:54*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[56*DATA_WIDTH-1:55*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[57*DATA_WIDTH-1:56*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[58*DATA_WIDTH-1:57*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[59*DATA_WIDTH-1:58*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[60*DATA_WIDTH-1:59*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[61*DATA_WIDTH-1:60*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[62*DATA_WIDTH-1:61*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[63*DATA_WIDTH-1:62*DATA_WIDTH] <= 0;
				reg_to_force_cache_LJ_Force_X[64*DATA_WIDTH-1:63*DATA_WIDTH] <= 0;
				reg_to_force_cache_particle_id[1*PARTICLE_ID_WIDTH-1:0*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[2*PARTICLE_ID_WIDTH-1:1*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[3*PARTICLE_ID_WIDTH-1:2*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[4*PARTICLE_ID_WIDTH-1:3*PARTICLE_ID_WIDTH] <= ref_particle_id_1_1;
				reg_to_force_cache_particle_id[5*PARTICLE_ID_WIDTH-1:4*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[6*PARTICLE_ID_WIDTH-1:5*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[7*PARTICLE_ID_WIDTH-1:6*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[8*PARTICLE_ID_WIDTH-1:7*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[9*PARTICLE_ID_WIDTH-1:8*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[10*PARTICLE_ID_WIDTH-1:9*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[11*PARTICLE_ID_WIDTH-1:10*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[12*PARTICLE_ID_WIDTH-1:11*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[13*PARTICLE_ID_WIDTH-1:12*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[14*PARTICLE_ID_WIDTH-1:13*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[15*PARTICLE_ID_WIDTH-1:14*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[16*PARTICLE_ID_WIDTH-1:15*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[17*PARTICLE_ID_WIDTH-1:16*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[18*PARTICLE_ID_WIDTH-1:17*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[19*PARTICLE_ID_WIDTH-1:18*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[20*PARTICLE_ID_WIDTH-1:19*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[21*PARTICLE_ID_WIDTH-1:20*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[22*PARTICLE_ID_WIDTH-1:21*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[23*PARTICLE_ID_WIDTH-1:22*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[24*PARTICLE_ID_WIDTH-1:23*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[25*PARTICLE_ID_WIDTH-1:24*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[26*PARTICLE_ID_WIDTH-1:25*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[27*PARTICLE_ID_WIDTH-1:26*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[28*PARTICLE_ID_WIDTH-1:27*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[29*PARTICLE_ID_WIDTH-1:28*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[30*PARTICLE_ID_WIDTH-1:29*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[31*PARTICLE_ID_WIDTH-1:30*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[32*PARTICLE_ID_WIDTH-1:31*PARTICLE_ID_WIDTH] <= neighbor_particle_id_1_1;
				reg_to_force_cache_particle_id[33*PARTICLE_ID_WIDTH-1:32*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[34*PARTICLE_ID_WIDTH-1:33*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[35*PARTICLE_ID_WIDTH-1:34*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[36*PARTICLE_ID_WIDTH-1:35*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[37*PARTICLE_ID_WIDTH-1:36*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[38*PARTICLE_ID_WIDTH-1:37*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[39*PARTICLE_ID_WIDTH-1:38*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[40*PARTICLE_ID_WIDTH-1:39*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[41*PARTICLE_ID_WIDTH-1:40*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[42*PARTICLE_ID_WIDTH-1:41*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[43*PARTICLE_ID_WIDTH-1:42*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[44*PARTICLE_ID_WIDTH-1:43*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[45*PARTICLE_ID_WIDTH-1:44*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[46*PARTICLE_ID_WIDTH-1:45*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[47*PARTICLE_ID_WIDTH-1:46*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[48*PARTICLE_ID_WIDTH-1:47*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[49*PARTICLE_ID_WIDTH-1:48*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[50*PARTICLE_ID_WIDTH-1:49*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[51*PARTICLE_ID_WIDTH-1:50*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[52*PARTICLE_ID_WIDTH-1:51*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[53*PARTICLE_ID_WIDTH-1:52*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[54*PARTICLE_ID_WIDTH-1:53*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[55*PARTICLE_ID_WIDTH-1:54*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[56*PARTICLE_ID_WIDTH-1:55*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[57*PARTICLE_ID_WIDTH-1:56*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[58*PARTICLE_ID_WIDTH-1:57*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[59*PARTICLE_ID_WIDTH-1:58*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[60*PARTICLE_ID_WIDTH-1:59*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[61*PARTICLE_ID_WIDTH-1:60*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[62*PARTICLE_ID_WIDTH-1:61*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[63*PARTICLE_ID_WIDTH-1:62*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_particle_id[64*PARTICLE_ID_WIDTH-1:63*PARTICLE_ID_WIDTH] <= 0;
				reg_to_force_cache_partial_force_valid[0] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[1] <= 1'b0;
				reg_to_force_cache_partial_force_valid[2] <= 1'b0;
				reg_to_force_cache_partial_force_valid[3] <= ref_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[4] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[5] <= 1'b0;
				reg_to_force_cache_partial_force_valid[6] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[7] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[8] <= 1'b0;
				reg_to_force_cache_partial_force_valid[9] <= 1'b0;
				reg_to_force_cache_partial_force_valid[10] <= 1'b0;
				reg_to_force_cache_partial_force_valid[11] <= 1'b0;
				reg_to_force_cache_partial_force_valid[12] <= 1'b0;
				reg_to_force_cache_partial_force_valid[13] <= 1'b0;
				reg_to_force_cache_partial_force_valid[14] <= 1'b0;
				reg_to_force_cache_partial_force_valid[15] <= 1'b0;
				reg_to_force_cache_partial_force_valid[16] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[17] <= 1'b0;
				reg_to_force_cache_partial_force_valid[18] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[19] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[20] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[21] <= 1'b0;
				reg_to_force_cache_partial_force_valid[22] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[23] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[24] <= 1'b0;
				reg_to_force_cache_partial_force_valid[25] <= 1'b0;
				reg_to_force_cache_partial_force_valid[26] <= 1'b0;
				reg_to_force_cache_partial_force_valid[27] <= 1'b0;
				reg_to_force_cache_partial_force_valid[28] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[29] <= 1'b0;
				reg_to_force_cache_partial_force_valid[30] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[31] <= neighbor_forceoutput_valid_1_1;
				reg_to_force_cache_partial_force_valid[32] <= 1'b0;
				reg_to_force_cache_partial_force_valid[33] <= 1'b0;
				reg_to_force_cache_partial_force_valid[34] <= 1'b0;
				reg_to_force_cache_partial_force_valid[35] <= 1'b0;
				reg_to_force_cache_partial_force_valid[36] <= 1'b0;
				reg_to_force_cache_partial_force_valid[37] <= 1'b0;
				reg_to_force_cache_partial_force_valid[38] <= 1'b0;
				reg_to_force_cache_partial_force_valid[39] <= 1'b0;
				reg_to_force_cache_partial_force_valid[40] <= 1'b0;
				reg_to_force_cache_partial_force_valid[41] <= 1'b0;
				reg_to_force_cache_partial_force_valid[42] <= 1'b0;
				reg_to_force_cache_partial_force_valid[43] <= 1'b0;
				reg_to_force_cache_partial_force_valid[44] <= 1'b0;
				reg_to_force_cache_partial_force_valid[45] <= 1'b0;
				reg_to_force_cache_partial_force_valid[46] <= 1'b0;
				reg_to_force_cache_partial_force_valid[47] <= 1'b0;
				reg_to_force_cache_partial_force_valid[48] <= 1'b0;
				reg_to_force_cache_partial_force_valid[49] <= 1'b0;
				reg_to_force_cache_partial_force_valid[50] <= 1'b0;
				reg_to_force_cache_partial_force_valid[51] <= 1'b0;
				reg_to_force_cache_partial_force_valid[52] <= 1'b0;
				reg_to_force_cache_partial_force_valid[53] <= 1'b0;
				reg_to_force_cache_partial_force_valid[54] <= 1'b0;
				reg_to_force_cache_partial_force_valid[55] <= 1'b0;
				reg_to_force_cache_partial_force_valid[56] <= 1'b0;
				reg_to_force_cache_partial_force_valid[57] <= 1'b0;
				reg_to_force_cache_partial_force_valid[58] <= 1'b0;
				reg_to_force_cache_partial_force_valid[59] <= 1'b0;
				reg_to_force_cache_partial_force_valid[60] <= 1'b0;
				reg_to_force_cache_partial_force_valid[61] <= 1'b0;
				reg_to_force_cache_partial_force_valid[62] <= 1'b0;
				reg_to_force_cache_partial_force_valid[63] <= 1'b0;
				reg_cells_to_pipeline_1_1 <= 	{
														Position_Cache_readout_position[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH],
														Position_Cache_readout_position[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH],
														Position_Cache_readout_position[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH],
														Position_Cache_readout_position[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH],
														Position_Cache_readout_position[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH],
														Position_Cache_readout_position[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH],
														Position_Cache_readout_position[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH],
														Position_Cache_readout_position[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH],
														Position_Cache_readout_position[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH],
														Position_Cache_readout_position[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH],
														Position_Cache_readout_position[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH],
														Position_Cache_readout_position[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH],
														Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH],
														Position_Cache_readout_position[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH]
														};
				reg_FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[2*CELL_ADDR_WIDTH-1:1*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[5*CELL_ADDR_WIDTH-1:4*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[3*CELL_ADDR_WIDTH-1:2*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[4*CELL_ADDR_WIDTH-1:3*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[15*CELL_ADDR_WIDTH-1:14*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[16*CELL_ADDR_WIDTH-1:15*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[17*CELL_ADDR_WIDTH-1:16*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[11*CELL_ADDR_WIDTH-1:10*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[18*CELL_ADDR_WIDTH-1:17*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[19*CELL_ADDR_WIDTH-1:18*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[9*CELL_ADDR_WIDTH-1:8*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[20*CELL_ADDR_WIDTH-1:19*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[10*CELL_ADDR_WIDTH-1:9*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[21*CELL_ADDR_WIDTH-1:20*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[14*CELL_ADDR_WIDTH-1:13*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[22*CELL_ADDR_WIDTH-1:21*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[23*CELL_ADDR_WIDTH-1:22*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[12*CELL_ADDR_WIDTH-1:11*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[24*CELL_ADDR_WIDTH-1:23*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[13*CELL_ADDR_WIDTH-1:12*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[25*CELL_ADDR_WIDTH-1:24*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[26*CELL_ADDR_WIDTH-1:25*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[27*CELL_ADDR_WIDTH-1:26*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[28*CELL_ADDR_WIDTH-1:27*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[29*CELL_ADDR_WIDTH-1:28*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[8*CELL_ADDR_WIDTH-1:7*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[30*CELL_ADDR_WIDTH-1:29*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[31*CELL_ADDR_WIDTH-1:30*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[6*CELL_ADDR_WIDTH-1:5*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[32*CELL_ADDR_WIDTH-1:31*CELL_ADDR_WIDTH] <= FSM_to_Cell_read_addr_1_1[7*CELL_ADDR_WIDTH-1:6*CELL_ADDR_WIDTH];
				reg_FSM_to_Cell_read_addr[33*CELL_ADDR_WIDTH-1:32*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[34*CELL_ADDR_WIDTH-1:33*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[35*CELL_ADDR_WIDTH-1:34*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[36*CELL_ADDR_WIDTH-1:35*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[37*CELL_ADDR_WIDTH-1:36*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[38*CELL_ADDR_WIDTH-1:37*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[39*CELL_ADDR_WIDTH-1:38*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[40*CELL_ADDR_WIDTH-1:39*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[41*CELL_ADDR_WIDTH-1:40*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[42*CELL_ADDR_WIDTH-1:41*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[43*CELL_ADDR_WIDTH-1:42*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[44*CELL_ADDR_WIDTH-1:43*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[45*CELL_ADDR_WIDTH-1:44*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[46*CELL_ADDR_WIDTH-1:45*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[47*CELL_ADDR_WIDTH-1:46*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[48*CELL_ADDR_WIDTH-1:47*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[49*CELL_ADDR_WIDTH-1:48*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[50*CELL_ADDR_WIDTH-1:49*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[51*CELL_ADDR_WIDTH-1:50*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[52*CELL_ADDR_WIDTH-1:51*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[53*CELL_ADDR_WIDTH-1:52*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[54*CELL_ADDR_WIDTH-1:53*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[55*CELL_ADDR_WIDTH-1:54*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[56*CELL_ADDR_WIDTH-1:55*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[57*CELL_ADDR_WIDTH-1:56*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[58*CELL_ADDR_WIDTH-1:57*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[59*CELL_ADDR_WIDTH-1:58*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[60*CELL_ADDR_WIDTH-1:59*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[61*CELL_ADDR_WIDTH-1:60*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[62*CELL_ADDR_WIDTH-1:61*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[63*CELL_ADDR_WIDTH-1:62*CELL_ADDR_WIDTH] <= 0;
				reg_FSM_to_Cell_read_addr[64*CELL_ADDR_WIDTH-1:63*CELL_ADDR_WIDTH] <= 0;
				if (FSM_to_Cell_rden_1_1)
					begin
					reg_FSM_to_Cell_rden[0] <= 1'b1;
					reg_FSM_to_Cell_rden[1] <= 1'b0;
					reg_FSM_to_Cell_rden[2] <= 1'b0;
					reg_FSM_to_Cell_rden[3] <= 1'b1;
					reg_FSM_to_Cell_rden[4] <= 1'b1;
					reg_FSM_to_Cell_rden[5] <= 1'b0;
					reg_FSM_to_Cell_rden[6] <= 1'b1;
					reg_FSM_to_Cell_rden[7] <= 1'b1;
					reg_FSM_to_Cell_rden[8] <= 1'b0;
					reg_FSM_to_Cell_rden[9] <= 1'b0;
					reg_FSM_to_Cell_rden[10] <= 1'b0;
					reg_FSM_to_Cell_rden[11] <= 1'b0;
					reg_FSM_to_Cell_rden[12] <= 1'b0;
					reg_FSM_to_Cell_rden[13] <= 1'b0;
					reg_FSM_to_Cell_rden[14] <= 1'b0;
					reg_FSM_to_Cell_rden[15] <= 1'b0;
					reg_FSM_to_Cell_rden[16] <= 1'b1;
					reg_FSM_to_Cell_rden[17] <= 1'b0;
					reg_FSM_to_Cell_rden[18] <= 1'b1;
					reg_FSM_to_Cell_rden[19] <= 1'b1;
					reg_FSM_to_Cell_rden[20] <= 1'b1;
					reg_FSM_to_Cell_rden[21] <= 1'b0;
					reg_FSM_to_Cell_rden[22] <= 1'b1;
					reg_FSM_to_Cell_rden[23] <= 1'b1;
					reg_FSM_to_Cell_rden[24] <= 1'b0;
					reg_FSM_to_Cell_rden[25] <= 1'b0;
					reg_FSM_to_Cell_rden[26] <= 1'b0;
					reg_FSM_to_Cell_rden[27] <= 1'b0;
					reg_FSM_to_Cell_rden[28] <= 1'b1;
					reg_FSM_to_Cell_rden[29] <= 1'b0;
					reg_FSM_to_Cell_rden[30] <= 1'b1;
					reg_FSM_to_Cell_rden[31] <= 1'b1;
					reg_FSM_to_Cell_rden[32] <= 1'b0;
					reg_FSM_to_Cell_rden[33] <= 1'b0;
					reg_FSM_to_Cell_rden[34] <= 1'b0;
					reg_FSM_to_Cell_rden[35] <= 1'b0;
					reg_FSM_to_Cell_rden[36] <= 1'b0;
					reg_FSM_to_Cell_rden[37] <= 1'b0;
					reg_FSM_to_Cell_rden[38] <= 1'b0;
					reg_FSM_to_Cell_rden[39] <= 1'b0;
					reg_FSM_to_Cell_rden[40] <= 1'b0;
					reg_FSM_to_Cell_rden[41] <= 1'b0;
					reg_FSM_to_Cell_rden[42] <= 1'b0;
					reg_FSM_to_Cell_rden[43] <= 1'b0;
					reg_FSM_to_Cell_rden[44] <= 1'b0;
					reg_FSM_to_Cell_rden[45] <= 1'b0;
					reg_FSM_to_Cell_rden[46] <= 1'b0;
					reg_FSM_to_Cell_rden[47] <= 1'b0;
					reg_FSM_to_Cell_rden[48] <= 1'b0;
					reg_FSM_to_Cell_rden[49] <= 1'b0;
					reg_FSM_to_Cell_rden[50] <= 1'b0;
					reg_FSM_to_Cell_rden[51] <= 1'b0;
					reg_FSM_to_Cell_rden[52] <= 1'b0;
					reg_FSM_to_Cell_rden[53] <= 1'b0;
					reg_FSM_to_Cell_rden[54] <= 1'b0;
					reg_FSM_to_Cell_rden[55] <= 1'b0;
					reg_FSM_to_Cell_rden[56] <= 1'b0;
					reg_FSM_to_Cell_rden[57] <= 1'b0;
					reg_FSM_to_Cell_rden[58] <= 1'b0;
					reg_FSM_to_Cell_rden[59] <= 1'b0;
					reg_FSM_to_Cell_rden[60] <= 1'b0;
					reg_FSM_to_Cell_rden[61] <= 1'b0;
					reg_FSM_to_Cell_rden[62] <= 1'b0;
					reg_FSM_to_Cell_rden[63] <= 1'b0;
					end
				else
					begin
					reg_FSM_to_Cell_rden[TOTAL_CELL_NUM-1:0] <= 0;
					end
				end
			default:
				begin
				reg_cells_to_pipeline_1_1 <= 0;
				reg_FSM_to_Cell_read_addr <= 0;
				reg_FSM_to_Cell_rden <= 0;
				reg_to_force_cache_partial_force_valid <= 0;
				reg_to_force_cache_particle_id <= 0;
				reg_to_force_cache_LJ_Force_Z <= 0;
				reg_to_force_cache_LJ_Force_Y <= 0;
				reg_to_force_cache_LJ_Force_X <= 0;
				end
			endcase
		end
	end
endmodule
