module TOP_RL_Pipeline_1st_Order
#(
	parameter DATA_WIDTH 				= 32,
	parameter INTERPOLATION_ORDER		= 1,
	parameter SEGMENT_NUM				= 12,
	parameter SEGMENT_WIDTH				= 4,
	parameter BIN_WIDTH					= 8,
	parameter BIN_NUM						= 256,
	parameter LOOKUP_NUM					= SEGMENT_NUM * BIN_NUM,			// SEGMENT_NUM * BIN_NUM
	parameter LOOKUP_ADDR_WIDTH		= SEGMENT_WIDTH + BIN_WIDTH		// log LOOKUP_NUM / log 2
)
(
	input  clk,
	input  rst,
	input  start,
	output [DATA_WIDTH-1:0] forceoutput,
	output forceoutput_valid,
	output done
);

	parameter PIPELINE_NUM = 200;

	wire [DATA_WIDTH-1:0] force_output_buffer [0:PIPELINE_NUM-1];
	wire [PIPELINE_NUM-1:0] force_valid;
	wire [PIPELINE_NUM-1:0] done_buffer;

	genvar i;
	for(i = 0; i < PIPELINE_NUM; i = i + 1)
	begin: generate_multiple_pipelines 
		RL_Pipeline_1st_Order
		#(
			DATA_WIDTH,
			INTERPOLATION_ORDER,
			SEGMENT_NUM,
			SEGMENT_WIDTH,
			BIN_WIDTH,
			BIN_NUM,
			LOOKUP_NUM,
			LOOKUP_ADDR_WIDTH
		)
		RL_Pipeline_1st_Order_inst
		(
			.clk(clk),
			.rst(rst),
			.start(start),
			.forceoutput(force_output_buffer[i]),
			.forceoutput_valid(force_valid[i]),
			.done(done_buffer[i])
		);
	end
	
	assign forceoutput = force_output_buffer[0] & force_output_buffer[1] & force_output_buffer[2] & force_output_buffer[3] & force_output_buffer[4] & force_output_buffer[5] & force_output_buffer[6] & force_output_buffer[7] & force_output_buffer[8] & force_output_buffer[9] & force_output_buffer[10] & force_output_buffer[11] & force_output_buffer[12] & force_output_buffer[13] & force_output_buffer[14] & force_output_buffer[15] & force_output_buffer[16] & force_output_buffer[17] & force_output_buffer[18] & force_output_buffer[19] & force_output_buffer[20] & force_output_buffer[21] & force_output_buffer[22] & force_output_buffer[23] & force_output_buffer[24] & force_output_buffer[25] & force_output_buffer[26] & force_output_buffer[27] & force_output_buffer[28] & force_output_buffer[29] & force_output_buffer[30] & force_output_buffer[31] & force_output_buffer[32] & force_output_buffer[33] & force_output_buffer[34] & force_output_buffer[35] & force_output_buffer[36] & force_output_buffer[37] & force_output_buffer[38] & force_output_buffer[39] & force_output_buffer[40] & force_output_buffer[41] & force_output_buffer[42] & force_output_buffer[43] & force_output_buffer[44] & force_output_buffer[45] & force_output_buffer[46] & force_output_buffer[47] & force_output_buffer[48] & force_output_buffer[49] & force_output_buffer[50] & force_output_buffer[51] & force_output_buffer[52] & force_output_buffer[53] & force_output_buffer[54] & force_output_buffer[55] & force_output_buffer[56] & force_output_buffer[57] & force_output_buffer[58] & force_output_buffer[59] & force_output_buffer[60] & force_output_buffer[61] & force_output_buffer[62] & force_output_buffer[63] & force_output_buffer[64] & force_output_buffer[65] & force_output_buffer[66] & force_output_buffer[67] & force_output_buffer[68] & force_output_buffer[69] & force_output_buffer[70] & force_output_buffer[71] & force_output_buffer[72] & force_output_buffer[73] & force_output_buffer[74] & force_output_buffer[75] & force_output_buffer[76] & force_output_buffer[77] & force_output_buffer[78] & force_output_buffer[79] & force_output_buffer[80] & force_output_buffer[81] & force_output_buffer[82] & force_output_buffer[83] & force_output_buffer[84] & force_output_buffer[85] & force_output_buffer[86] & force_output_buffer[87] & force_output_buffer[88] & force_output_buffer[89] & force_output_buffer[90] & force_output_buffer[91] & force_output_buffer[92] & force_output_buffer[93] & force_output_buffer[94] & force_output_buffer[95] & force_output_buffer[96] & force_output_buffer[97] & force_output_buffer[98] & force_output_buffer[99] & force_output_buffer[100] & force_output_buffer[101] & force_output_buffer[102] & force_output_buffer[103] & force_output_buffer[104] & force_output_buffer[105] & force_output_buffer[106] & force_output_buffer[107] & force_output_buffer[108] & force_output_buffer[109] & force_output_buffer[110] & force_output_buffer[111] & force_output_buffer[112] & force_output_buffer[113] & force_output_buffer[114] & force_output_buffer[115] & force_output_buffer[116] & force_output_buffer[117] & force_output_buffer[118] & force_output_buffer[119] & force_output_buffer[120] & force_output_buffer[121] & force_output_buffer[122] & force_output_buffer[123] & force_output_buffer[124] & force_output_buffer[125] & force_output_buffer[126] & force_output_buffer[127] & force_output_buffer[128] & force_output_buffer[129] & force_output_buffer[130] & force_output_buffer[131] & force_output_buffer[132] & force_output_buffer[133] & force_output_buffer[134] & force_output_buffer[135] & force_output_buffer[136] & force_output_buffer[137] & force_output_buffer[138] & force_output_buffer[139] & force_output_buffer[140] & force_output_buffer[141] & force_output_buffer[142] & force_output_buffer[143] & force_output_buffer[144] & force_output_buffer[145] & force_output_buffer[146] & force_output_buffer[147] & force_output_buffer[148] & force_output_buffer[149] & force_output_buffer[150] & force_output_buffer[151] & force_output_buffer[152] & force_output_buffer[153] & force_output_buffer[154] & force_output_buffer[155] & force_output_buffer[156] & force_output_buffer[157] & force_output_buffer[158] & force_output_buffer[159] & force_output_buffer[160] & force_output_buffer[161] & force_output_buffer[162] & force_output_buffer[163] & force_output_buffer[164] & force_output_buffer[165] & force_output_buffer[166] & force_output_buffer[167] & force_output_buffer[168] & force_output_buffer[169] & force_output_buffer[170] & force_output_buffer[171] & force_output_buffer[172] & force_output_buffer[173] & force_output_buffer[174] & force_output_buffer[175] & force_output_buffer[176] & force_output_buffer[177] & force_output_buffer[178] & force_output_buffer[179] & force_output_buffer[180] & force_output_buffer[181] & force_output_buffer[182] & force_output_buffer[183] & force_output_buffer[184] & force_output_buffer[185] & force_output_buffer[186] & force_output_buffer[187] & force_output_buffer[188] & force_output_buffer[189] & force_output_buffer[190] & force_output_buffer[191] & force_output_buffer[192] & force_output_buffer[193] & force_output_buffer[194] & force_output_buffer[195] & force_output_buffer[196] & force_output_buffer[197] & force_output_buffer[198] & force_output_buffer[199];
	assign forceoutput_valid = force_output_buffer[0] & force_output_buffer[1] & force_output_buffer[2] & force_output_buffer[3] & force_output_buffer[4] & force_output_buffer[5] & force_output_buffer[6] & force_output_buffer[7] & force_output_buffer[8] & force_output_buffer[9] & force_output_buffer[10] & force_output_buffer[11] & force_output_buffer[12] & force_output_buffer[13] & force_output_buffer[14] & force_output_buffer[15] & force_output_buffer[16] & force_output_buffer[17] & force_output_buffer[18] & force_output_buffer[19] & force_output_buffer[20] & force_output_buffer[21] & force_output_buffer[22] & force_output_buffer[23] & force_output_buffer[24] & force_output_buffer[25] & force_output_buffer[26] & force_output_buffer[27] & force_output_buffer[28] & force_output_buffer[29] & force_output_buffer[30] & force_output_buffer[31] & force_output_buffer[32] & force_output_buffer[33] & force_output_buffer[34] & force_output_buffer[35] & force_output_buffer[36] & force_output_buffer[37] & force_output_buffer[38] & force_output_buffer[39] & force_output_buffer[40] & force_output_buffer[41] & force_output_buffer[42] & force_output_buffer[43] & force_output_buffer[44] & force_output_buffer[45] & force_output_buffer[46] & force_output_buffer[47] & force_output_buffer[48] & force_output_buffer[49] & force_output_buffer[50] & force_output_buffer[51] & force_output_buffer[52] & force_output_buffer[53] & force_output_buffer[54] & force_output_buffer[55] & force_output_buffer[56] & force_output_buffer[57] & force_output_buffer[58] & force_output_buffer[59] & force_output_buffer[60] & force_output_buffer[61] & force_output_buffer[62] & force_output_buffer[63] & force_output_buffer[64] & force_output_buffer[65] & force_output_buffer[66] & force_output_buffer[67] & force_output_buffer[68] & force_output_buffer[69] & force_output_buffer[70] & force_output_buffer[71] & force_output_buffer[72] & force_output_buffer[73] & force_output_buffer[74] & force_output_buffer[75] & force_output_buffer[76] & force_output_buffer[77] & force_output_buffer[78] & force_output_buffer[79] & force_output_buffer[80] & force_output_buffer[81] & force_output_buffer[82] & force_output_buffer[83] & force_output_buffer[84] & force_output_buffer[85] & force_output_buffer[86] & force_output_buffer[87] & force_output_buffer[88] & force_output_buffer[89] & force_output_buffer[90] & force_output_buffer[91] & force_output_buffer[92] & force_output_buffer[93] & force_output_buffer[94] & force_output_buffer[95] & force_output_buffer[96] & force_output_buffer[97] & force_output_buffer[98] & force_output_buffer[99] & force_output_buffer[100] & force_output_buffer[101] & force_output_buffer[102] & force_output_buffer[103] & force_output_buffer[104] & force_output_buffer[105] & force_output_buffer[106] & force_output_buffer[107] & force_output_buffer[108] & force_output_buffer[109] & force_output_buffer[110] & force_output_buffer[111] & force_output_buffer[112] & force_output_buffer[113] & force_output_buffer[114] & force_output_buffer[115] & force_output_buffer[116] & force_output_buffer[117] & force_output_buffer[118] & force_output_buffer[119] & force_output_buffer[120] & force_output_buffer[121] & force_output_buffer[122] & force_output_buffer[123] & force_output_buffer[124] & force_output_buffer[125] & force_output_buffer[126] & force_output_buffer[127] & force_output_buffer[128] & force_output_buffer[129] & force_output_buffer[130] & force_output_buffer[131] & force_output_buffer[132] & force_output_buffer[133] & force_output_buffer[134] & force_output_buffer[135] & force_output_buffer[136] & force_output_buffer[137] & force_output_buffer[138] & force_output_buffer[139] & force_output_buffer[140] & force_output_buffer[141] & force_output_buffer[142] & force_output_buffer[143] & force_output_buffer[144] & force_output_buffer[145] & force_output_buffer[146] & force_output_buffer[147] & force_output_buffer[148] & force_output_buffer[149] & force_output_buffer[150] & force_output_buffer[151] & force_output_buffer[152] & force_output_buffer[153] & force_output_buffer[154] & force_output_buffer[155] & force_output_buffer[156] & force_output_buffer[157] & force_output_buffer[158] & force_output_buffer[159] & force_output_buffer[160] & force_output_buffer[161] & force_output_buffer[162] & force_output_buffer[163] & force_output_buffer[164] & force_output_buffer[165] & force_output_buffer[166] & force_output_buffer[167] & force_output_buffer[168] & force_output_buffer[169] & force_output_buffer[170] & force_output_buffer[171] & force_output_buffer[172] & force_output_buffer[173] & force_output_buffer[174] & force_output_buffer[175] & force_output_buffer[176] & force_output_buffer[177] & force_output_buffer[178] & force_output_buffer[179] & force_output_buffer[180] & force_output_buffer[181] & force_output_buffer[182] & force_output_buffer[183] & force_output_buffer[184] & force_output_buffer[185] & force_output_buffer[186] & force_output_buffer[187] & force_output_buffer[188] & force_output_buffer[189] & force_output_buffer[190] & force_output_buffer[191] & force_output_buffer[192] & force_output_buffer[193] & force_output_buffer[194] & force_output_buffer[195] & force_output_buffer[196] & force_output_buffer[197] & force_output_buffer[198] & force_output_buffer[199];
	assign done = done_buffer[0] & done_buffer[1] & done_buffer[2] & done_buffer[3] & done_buffer[4] & done_buffer[5] & done_buffer[6] & done_buffer[7] & done_buffer[8] & done_buffer[9] & done_buffer[10] & done_buffer[11] & done_buffer[12] & done_buffer[13] & done_buffer[14] & done_buffer[15] & done_buffer[16] & done_buffer[17] & done_buffer[18] & done_buffer[19] & done_buffer[20] & done_buffer[21] & done_buffer[22] & done_buffer[23] & done_buffer[24] & done_buffer[25] & done_buffer[26] & done_buffer[27] & done_buffer[28] & done_buffer[29] & done_buffer[30] & done_buffer[31] & done_buffer[32] & done_buffer[33] & done_buffer[34] & done_buffer[35] & done_buffer[36] & done_buffer[37] & done_buffer[38] & done_buffer[39] & done_buffer[40] & done_buffer[41] & done_buffer[42] & done_buffer[43] & done_buffer[44] & done_buffer[45] & done_buffer[46] & done_buffer[47] & done_buffer[48] & done_buffer[49] & done_buffer[50] & done_buffer[51] & done_buffer[52] & done_buffer[53] & done_buffer[54] & done_buffer[55] & done_buffer[56] & done_buffer[57] & done_buffer[58] & done_buffer[59] & done_buffer[60] & done_buffer[61] & done_buffer[62] & done_buffer[63] & done_buffer[64] & done_buffer[65] & done_buffer[66] & done_buffer[67] & done_buffer[68] & done_buffer[69] & done_buffer[70] & done_buffer[71] & done_buffer[72] & done_buffer[73] & done_buffer[74] & done_buffer[75] & done_buffer[76] & done_buffer[77] & done_buffer[78] & done_buffer[79] & done_buffer[80] & done_buffer[81] & done_buffer[82] & done_buffer[83] & done_buffer[84] & done_buffer[85] & done_buffer[86] & done_buffer[87] & done_buffer[88] & done_buffer[89] & done_buffer[90] & done_buffer[91] & done_buffer[92] & done_buffer[93] & done_buffer[94] & done_buffer[95] & done_buffer[96] & done_buffer[97] & done_buffer[98] & done_buffer[99] & done_buffer[100] & done_buffer[101] & done_buffer[102] & done_buffer[103] & done_buffer[104] & done_buffer[105] & done_buffer[106] & done_buffer[107] & done_buffer[108] & done_buffer[109] & done_buffer[110] & done_buffer[111] & done_buffer[112] & done_buffer[113] & done_buffer[114] & done_buffer[115] & done_buffer[116] & done_buffer[117] & done_buffer[118] & done_buffer[119] & done_buffer[120] & done_buffer[121] & done_buffer[122] & done_buffer[123] & done_buffer[124] & done_buffer[125] & done_buffer[126] & done_buffer[127] & done_buffer[128] & done_buffer[129] & done_buffer[130] & done_buffer[131] & done_buffer[132] & done_buffer[133] & done_buffer[134] & done_buffer[135] & done_buffer[136] & done_buffer[137] & done_buffer[138] & done_buffer[139] & done_buffer[140] & done_buffer[141] & done_buffer[142] & done_buffer[143] & done_buffer[144] & done_buffer[145] & done_buffer[146] & done_buffer[147] & done_buffer[148] & done_buffer[149] & done_buffer[150] & done_buffer[151] & done_buffer[152] & done_buffer[153] & done_buffer[154] & done_buffer[155] & done_buffer[156] & done_buffer[157] & done_buffer[158] & done_buffer[159] & done_buffer[160] & done_buffer[161] & done_buffer[162] & done_buffer[163] & done_buffer[164] & done_buffer[165] & done_buffer[166] & done_buffer[167] & done_buffer[168] & done_buffer[169] & done_buffer[170] & done_buffer[171] & done_buffer[172] & done_buffer[173] & done_buffer[174] & done_buffer[175] & done_buffer[176] & done_buffer[177] & done_buffer[178] & done_buffer[179] & done_buffer[180] & done_buffer[181] & done_buffer[182] & done_buffer[183] & done_buffer[184] & done_buffer[185] & done_buffer[186] & done_buffer[187] & done_buffer[188] & done_buffer[189] & done_buffer[190] & done_buffer[191] & done_buffer[192] & done_buffer[193] & done_buffer[194] & done_buffer[195] & done_buffer[196] & done_buffer[197] & done_buffer[198] & done_buffer[199];
endmodule