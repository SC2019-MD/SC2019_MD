/*****************************************************
Used to store all the force caches, nice and clean
*****************************************************/


module All_Force_Caches_64_Cells
#(
	parameter DATA_WIDTH 					= 32,
	parameter TOTAL_CELL_NUM				= 64,
	parameter FORCE_CACHE_BUFFER_DEPTH	= 16,
	parameter FORCE_CACHE_BUFFER_ADDR_WIDTH = 4,	
	parameter CELL_ID_WIDTH					= 4,
	parameter MAX_CELL_PARTICLE_NUM		= 290,
	parameter CELL_ADDR_WIDTH				= 9,
	parameter PARTICLE_ID_WIDTH			= CELL_ID_WIDTH*3+CELL_ADDR_WIDTH, 
	
	parameter FORCE_EVAL_FIFO_DATA_WIDTH = 113
)
(
	input clk, 
	input rst, 
	input [TOTAL_CELL_NUM-1:0] wire_motion_update_to_cache_read_force_request,
	input [CELL_ADDR_WIDTH-1:0]Motion_Update_force_read_addr,
	input [TOTAL_CELL_NUM*FORCE_EVAL_FIFO_DATA_WIDTH-1:0] valid_force_values,
	
	output [TOTAL_CELL_NUM*3*DATA_WIDTH-1:0] wire_cache_to_motion_update_partial_force,
	output [TOTAL_CELL_NUM*PARTICLE_ID_WIDTH-1:0] wire_cache_to_motion_update_particle_id,
	output [TOTAL_CELL_NUM-1:0] wire_cache_to_motion_update_partial_force_valid
);
	
	wire [TOTAL_CELL_NUM*DATA_WIDTH-1:0] to_force_cache_LJ_Force_Z;
	wire [TOTAL_CELL_NUM*DATA_WIDTH-1:0] to_force_cache_LJ_Force_Y;
	wire [TOTAL_CELL_NUM*DATA_WIDTH-1:0] to_force_cache_LJ_Force_X;
	wire [TOTAL_CELL_NUM-1:0] to_force_cache_partial_force_valid;
	wire [TOTAL_CELL_NUM*PARTICLE_ID_WIDTH-1:0] to_force_cache_particle_id;
	
	assign to_force_cache_LJ_Force_Z[1*DATA_WIDTH-1:0*DATA_WIDTH] = valid_force_values[1*FORCE_EVAL_FIFO_DATA_WIDTH-1:0*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[2*DATA_WIDTH-1:1*DATA_WIDTH] = valid_force_values[2*FORCE_EVAL_FIFO_DATA_WIDTH-1:1*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[3*DATA_WIDTH-1:2*DATA_WIDTH] = valid_force_values[3*FORCE_EVAL_FIFO_DATA_WIDTH-1:2*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[4*DATA_WIDTH-1:3*DATA_WIDTH] = valid_force_values[4*FORCE_EVAL_FIFO_DATA_WIDTH-1:3*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[5*DATA_WIDTH-1:4*DATA_WIDTH] = valid_force_values[5*FORCE_EVAL_FIFO_DATA_WIDTH-1:4*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[6*DATA_WIDTH-1:5*DATA_WIDTH] = valid_force_values[6*FORCE_EVAL_FIFO_DATA_WIDTH-1:5*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[7*DATA_WIDTH-1:6*DATA_WIDTH] = valid_force_values[7*FORCE_EVAL_FIFO_DATA_WIDTH-1:6*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[8*DATA_WIDTH-1:7*DATA_WIDTH] = valid_force_values[8*FORCE_EVAL_FIFO_DATA_WIDTH-1:7*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[9*DATA_WIDTH-1:8*DATA_WIDTH] = valid_force_values[9*FORCE_EVAL_FIFO_DATA_WIDTH-1:8*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[10*DATA_WIDTH-1:9*DATA_WIDTH] = valid_force_values[10*FORCE_EVAL_FIFO_DATA_WIDTH-1:9*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[11*DATA_WIDTH-1:10*DATA_WIDTH] = valid_force_values[11*FORCE_EVAL_FIFO_DATA_WIDTH-1:10*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[12*DATA_WIDTH-1:11*DATA_WIDTH] = valid_force_values[12*FORCE_EVAL_FIFO_DATA_WIDTH-1:11*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[13*DATA_WIDTH-1:12*DATA_WIDTH] = valid_force_values[13*FORCE_EVAL_FIFO_DATA_WIDTH-1:12*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[14*DATA_WIDTH-1:13*DATA_WIDTH] = valid_force_values[14*FORCE_EVAL_FIFO_DATA_WIDTH-1:13*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[15*DATA_WIDTH-1:14*DATA_WIDTH] = valid_force_values[15*FORCE_EVAL_FIFO_DATA_WIDTH-1:14*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[16*DATA_WIDTH-1:15*DATA_WIDTH] = valid_force_values[16*FORCE_EVAL_FIFO_DATA_WIDTH-1:15*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[17*DATA_WIDTH-1:16*DATA_WIDTH] = valid_force_values[17*FORCE_EVAL_FIFO_DATA_WIDTH-1:16*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[18*DATA_WIDTH-1:17*DATA_WIDTH] = valid_force_values[18*FORCE_EVAL_FIFO_DATA_WIDTH-1:17*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[19*DATA_WIDTH-1:18*DATA_WIDTH] = valid_force_values[19*FORCE_EVAL_FIFO_DATA_WIDTH-1:18*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[20*DATA_WIDTH-1:19*DATA_WIDTH] = valid_force_values[20*FORCE_EVAL_FIFO_DATA_WIDTH-1:19*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[21*DATA_WIDTH-1:20*DATA_WIDTH] = valid_force_values[21*FORCE_EVAL_FIFO_DATA_WIDTH-1:20*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[22*DATA_WIDTH-1:21*DATA_WIDTH] = valid_force_values[22*FORCE_EVAL_FIFO_DATA_WIDTH-1:21*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[23*DATA_WIDTH-1:22*DATA_WIDTH] = valid_force_values[23*FORCE_EVAL_FIFO_DATA_WIDTH-1:22*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[24*DATA_WIDTH-1:23*DATA_WIDTH] = valid_force_values[24*FORCE_EVAL_FIFO_DATA_WIDTH-1:23*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[25*DATA_WIDTH-1:24*DATA_WIDTH] = valid_force_values[25*FORCE_EVAL_FIFO_DATA_WIDTH-1:24*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[26*DATA_WIDTH-1:25*DATA_WIDTH] = valid_force_values[26*FORCE_EVAL_FIFO_DATA_WIDTH-1:25*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[27*DATA_WIDTH-1:26*DATA_WIDTH] = valid_force_values[27*FORCE_EVAL_FIFO_DATA_WIDTH-1:26*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[28*DATA_WIDTH-1:27*DATA_WIDTH] = valid_force_values[28*FORCE_EVAL_FIFO_DATA_WIDTH-1:27*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[29*DATA_WIDTH-1:28*DATA_WIDTH] = valid_force_values[29*FORCE_EVAL_FIFO_DATA_WIDTH-1:28*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[30*DATA_WIDTH-1:29*DATA_WIDTH] = valid_force_values[30*FORCE_EVAL_FIFO_DATA_WIDTH-1:29*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[31*DATA_WIDTH-1:30*DATA_WIDTH] = valid_force_values[31*FORCE_EVAL_FIFO_DATA_WIDTH-1:30*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[32*DATA_WIDTH-1:31*DATA_WIDTH] = valid_force_values[32*FORCE_EVAL_FIFO_DATA_WIDTH-1:31*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[33*DATA_WIDTH-1:32*DATA_WIDTH] = valid_force_values[33*FORCE_EVAL_FIFO_DATA_WIDTH-1:32*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[34*DATA_WIDTH-1:33*DATA_WIDTH] = valid_force_values[34*FORCE_EVAL_FIFO_DATA_WIDTH-1:33*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[35*DATA_WIDTH-1:34*DATA_WIDTH] = valid_force_values[35*FORCE_EVAL_FIFO_DATA_WIDTH-1:34*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[36*DATA_WIDTH-1:35*DATA_WIDTH] = valid_force_values[36*FORCE_EVAL_FIFO_DATA_WIDTH-1:35*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[37*DATA_WIDTH-1:36*DATA_WIDTH] = valid_force_values[37*FORCE_EVAL_FIFO_DATA_WIDTH-1:36*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[38*DATA_WIDTH-1:37*DATA_WIDTH] = valid_force_values[38*FORCE_EVAL_FIFO_DATA_WIDTH-1:37*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[39*DATA_WIDTH-1:38*DATA_WIDTH] = valid_force_values[39*FORCE_EVAL_FIFO_DATA_WIDTH-1:38*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[40*DATA_WIDTH-1:39*DATA_WIDTH] = valid_force_values[40*FORCE_EVAL_FIFO_DATA_WIDTH-1:39*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[41*DATA_WIDTH-1:40*DATA_WIDTH] = valid_force_values[41*FORCE_EVAL_FIFO_DATA_WIDTH-1:40*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[42*DATA_WIDTH-1:41*DATA_WIDTH] = valid_force_values[42*FORCE_EVAL_FIFO_DATA_WIDTH-1:41*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[43*DATA_WIDTH-1:42*DATA_WIDTH] = valid_force_values[43*FORCE_EVAL_FIFO_DATA_WIDTH-1:42*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[44*DATA_WIDTH-1:43*DATA_WIDTH] = valid_force_values[44*FORCE_EVAL_FIFO_DATA_WIDTH-1:43*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[45*DATA_WIDTH-1:44*DATA_WIDTH] = valid_force_values[45*FORCE_EVAL_FIFO_DATA_WIDTH-1:44*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[46*DATA_WIDTH-1:45*DATA_WIDTH] = valid_force_values[46*FORCE_EVAL_FIFO_DATA_WIDTH-1:45*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[47*DATA_WIDTH-1:46*DATA_WIDTH] = valid_force_values[47*FORCE_EVAL_FIFO_DATA_WIDTH-1:46*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[48*DATA_WIDTH-1:47*DATA_WIDTH] = valid_force_values[48*FORCE_EVAL_FIFO_DATA_WIDTH-1:47*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[49*DATA_WIDTH-1:48*DATA_WIDTH] = valid_force_values[49*FORCE_EVAL_FIFO_DATA_WIDTH-1:48*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[50*DATA_WIDTH-1:49*DATA_WIDTH] = valid_force_values[50*FORCE_EVAL_FIFO_DATA_WIDTH-1:49*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[51*DATA_WIDTH-1:50*DATA_WIDTH] = valid_force_values[51*FORCE_EVAL_FIFO_DATA_WIDTH-1:50*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[52*DATA_WIDTH-1:51*DATA_WIDTH] = valid_force_values[52*FORCE_EVAL_FIFO_DATA_WIDTH-1:51*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[53*DATA_WIDTH-1:52*DATA_WIDTH] = valid_force_values[53*FORCE_EVAL_FIFO_DATA_WIDTH-1:52*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[54*DATA_WIDTH-1:53*DATA_WIDTH] = valid_force_values[54*FORCE_EVAL_FIFO_DATA_WIDTH-1:53*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[55*DATA_WIDTH-1:54*DATA_WIDTH] = valid_force_values[55*FORCE_EVAL_FIFO_DATA_WIDTH-1:54*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[56*DATA_WIDTH-1:55*DATA_WIDTH] = valid_force_values[56*FORCE_EVAL_FIFO_DATA_WIDTH-1:55*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[57*DATA_WIDTH-1:56*DATA_WIDTH] = valid_force_values[57*FORCE_EVAL_FIFO_DATA_WIDTH-1:56*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[58*DATA_WIDTH-1:57*DATA_WIDTH] = valid_force_values[58*FORCE_EVAL_FIFO_DATA_WIDTH-1:57*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[59*DATA_WIDTH-1:58*DATA_WIDTH] = valid_force_values[59*FORCE_EVAL_FIFO_DATA_WIDTH-1:58*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[60*DATA_WIDTH-1:59*DATA_WIDTH] = valid_force_values[60*FORCE_EVAL_FIFO_DATA_WIDTH-1:59*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[61*DATA_WIDTH-1:60*DATA_WIDTH] = valid_force_values[61*FORCE_EVAL_FIFO_DATA_WIDTH-1:60*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[62*DATA_WIDTH-1:61*DATA_WIDTH] = valid_force_values[62*FORCE_EVAL_FIFO_DATA_WIDTH-1:61*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[63*DATA_WIDTH-1:62*DATA_WIDTH] = valid_force_values[63*FORCE_EVAL_FIFO_DATA_WIDTH-1:62*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Z[64*DATA_WIDTH-1:63*DATA_WIDTH] = valid_force_values[64*FORCE_EVAL_FIFO_DATA_WIDTH-1:63*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+2*DATA_WIDTH+1];

	assign to_force_cache_LJ_Force_Y[1*DATA_WIDTH-1:0*DATA_WIDTH] = valid_force_values[1*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:0*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[2*DATA_WIDTH-1:1*DATA_WIDTH] = valid_force_values[2*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:1*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[3*DATA_WIDTH-1:2*DATA_WIDTH] = valid_force_values[3*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:2*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[4*DATA_WIDTH-1:3*DATA_WIDTH] = valid_force_values[4*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:3*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[5*DATA_WIDTH-1:4*DATA_WIDTH] = valid_force_values[5*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:4*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[6*DATA_WIDTH-1:5*DATA_WIDTH] = valid_force_values[6*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:5*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[7*DATA_WIDTH-1:6*DATA_WIDTH] = valid_force_values[7*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:6*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[8*DATA_WIDTH-1:7*DATA_WIDTH] = valid_force_values[8*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:7*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[9*DATA_WIDTH-1:8*DATA_WIDTH] = valid_force_values[9*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:8*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[10*DATA_WIDTH-1:9*DATA_WIDTH] = valid_force_values[10*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:9*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[11*DATA_WIDTH-1:10*DATA_WIDTH] = valid_force_values[11*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:10*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[12*DATA_WIDTH-1:11*DATA_WIDTH] = valid_force_values[12*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:11*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[13*DATA_WIDTH-1:12*DATA_WIDTH] = valid_force_values[13*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:12*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[14*DATA_WIDTH-1:13*DATA_WIDTH] = valid_force_values[14*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:13*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[15*DATA_WIDTH-1:14*DATA_WIDTH] = valid_force_values[15*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:14*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[16*DATA_WIDTH-1:15*DATA_WIDTH] = valid_force_values[16*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:15*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[17*DATA_WIDTH-1:16*DATA_WIDTH] = valid_force_values[17*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:16*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[18*DATA_WIDTH-1:17*DATA_WIDTH] = valid_force_values[18*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:17*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[19*DATA_WIDTH-1:18*DATA_WIDTH] = valid_force_values[19*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:18*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[20*DATA_WIDTH-1:19*DATA_WIDTH] = valid_force_values[20*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:19*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[21*DATA_WIDTH-1:20*DATA_WIDTH] = valid_force_values[21*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:20*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[22*DATA_WIDTH-1:21*DATA_WIDTH] = valid_force_values[22*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:21*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[23*DATA_WIDTH-1:22*DATA_WIDTH] = valid_force_values[23*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:22*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[24*DATA_WIDTH-1:23*DATA_WIDTH] = valid_force_values[24*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:23*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[25*DATA_WIDTH-1:24*DATA_WIDTH] = valid_force_values[25*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:24*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[26*DATA_WIDTH-1:25*DATA_WIDTH] = valid_force_values[26*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:25*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[27*DATA_WIDTH-1:26*DATA_WIDTH] = valid_force_values[27*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:26*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[28*DATA_WIDTH-1:27*DATA_WIDTH] = valid_force_values[28*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:27*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[29*DATA_WIDTH-1:28*DATA_WIDTH] = valid_force_values[29*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:28*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[30*DATA_WIDTH-1:29*DATA_WIDTH] = valid_force_values[30*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:29*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[31*DATA_WIDTH-1:30*DATA_WIDTH] = valid_force_values[31*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:30*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[32*DATA_WIDTH-1:31*DATA_WIDTH] = valid_force_values[32*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:31*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[33*DATA_WIDTH-1:32*DATA_WIDTH] = valid_force_values[33*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:32*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[34*DATA_WIDTH-1:33*DATA_WIDTH] = valid_force_values[34*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:33*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[35*DATA_WIDTH-1:34*DATA_WIDTH] = valid_force_values[35*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:34*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[36*DATA_WIDTH-1:35*DATA_WIDTH] = valid_force_values[36*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:35*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[37*DATA_WIDTH-1:36*DATA_WIDTH] = valid_force_values[37*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:36*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[38*DATA_WIDTH-1:37*DATA_WIDTH] = valid_force_values[38*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:37*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[39*DATA_WIDTH-1:38*DATA_WIDTH] = valid_force_values[39*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:38*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[40*DATA_WIDTH-1:39*DATA_WIDTH] = valid_force_values[40*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:39*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[41*DATA_WIDTH-1:40*DATA_WIDTH] = valid_force_values[41*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:40*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[42*DATA_WIDTH-1:41*DATA_WIDTH] = valid_force_values[42*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:41*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[43*DATA_WIDTH-1:42*DATA_WIDTH] = valid_force_values[43*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:42*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[44*DATA_WIDTH-1:43*DATA_WIDTH] = valid_force_values[44*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:43*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[45*DATA_WIDTH-1:44*DATA_WIDTH] = valid_force_values[45*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:44*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[46*DATA_WIDTH-1:45*DATA_WIDTH] = valid_force_values[46*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:45*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[47*DATA_WIDTH-1:46*DATA_WIDTH] = valid_force_values[47*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:46*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[48*DATA_WIDTH-1:47*DATA_WIDTH] = valid_force_values[48*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:47*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[49*DATA_WIDTH-1:48*DATA_WIDTH] = valid_force_values[49*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:48*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[50*DATA_WIDTH-1:49*DATA_WIDTH] = valid_force_values[50*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:49*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[51*DATA_WIDTH-1:50*DATA_WIDTH] = valid_force_values[51*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:50*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[52*DATA_WIDTH-1:51*DATA_WIDTH] = valid_force_values[52*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:51*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[53*DATA_WIDTH-1:52*DATA_WIDTH] = valid_force_values[53*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:52*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[54*DATA_WIDTH-1:53*DATA_WIDTH] = valid_force_values[54*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:53*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[55*DATA_WIDTH-1:54*DATA_WIDTH] = valid_force_values[55*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:54*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[56*DATA_WIDTH-1:55*DATA_WIDTH] = valid_force_values[56*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:55*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[57*DATA_WIDTH-1:56*DATA_WIDTH] = valid_force_values[57*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:56*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[58*DATA_WIDTH-1:57*DATA_WIDTH] = valid_force_values[58*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:57*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[59*DATA_WIDTH-1:58*DATA_WIDTH] = valid_force_values[59*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:58*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[60*DATA_WIDTH-1:59*DATA_WIDTH] = valid_force_values[60*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:59*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[61*DATA_WIDTH-1:60*DATA_WIDTH] = valid_force_values[61*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:60*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[62*DATA_WIDTH-1:61*DATA_WIDTH] = valid_force_values[62*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:61*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[63*DATA_WIDTH-1:62*DATA_WIDTH] = valid_force_values[63*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:62*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	assign to_force_cache_LJ_Force_Y[64*DATA_WIDTH-1:63*DATA_WIDTH] = valid_force_values[64*FORCE_EVAL_FIFO_DATA_WIDTH-DATA_WIDTH-1:63*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+DATA_WIDTH+1];
	
	assign to_force_cache_LJ_Force_X[1*DATA_WIDTH-1:0*DATA_WIDTH] = valid_force_values[1*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:0*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[2*DATA_WIDTH-1:1*DATA_WIDTH] = valid_force_values[2*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:1*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[3*DATA_WIDTH-1:2*DATA_WIDTH] = valid_force_values[3*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:2*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[4*DATA_WIDTH-1:3*DATA_WIDTH] = valid_force_values[4*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:3*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[5*DATA_WIDTH-1:4*DATA_WIDTH] = valid_force_values[5*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:4*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[6*DATA_WIDTH-1:5*DATA_WIDTH] = valid_force_values[6*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:5*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[7*DATA_WIDTH-1:6*DATA_WIDTH] = valid_force_values[7*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:6*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[8*DATA_WIDTH-1:7*DATA_WIDTH] = valid_force_values[8*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:7*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[9*DATA_WIDTH-1:8*DATA_WIDTH] = valid_force_values[9*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:8*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[10*DATA_WIDTH-1:9*DATA_WIDTH] = valid_force_values[10*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:9*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[11*DATA_WIDTH-1:10*DATA_WIDTH] = valid_force_values[11*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:10*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[12*DATA_WIDTH-1:11*DATA_WIDTH] = valid_force_values[12*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:11*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[13*DATA_WIDTH-1:12*DATA_WIDTH] = valid_force_values[13*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:12*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[14*DATA_WIDTH-1:13*DATA_WIDTH] = valid_force_values[14*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:13*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[15*DATA_WIDTH-1:14*DATA_WIDTH] = valid_force_values[15*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:14*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[16*DATA_WIDTH-1:15*DATA_WIDTH] = valid_force_values[16*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:15*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[17*DATA_WIDTH-1:16*DATA_WIDTH] = valid_force_values[17*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:16*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[18*DATA_WIDTH-1:17*DATA_WIDTH] = valid_force_values[18*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:17*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[19*DATA_WIDTH-1:18*DATA_WIDTH] = valid_force_values[19*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:18*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[20*DATA_WIDTH-1:19*DATA_WIDTH] = valid_force_values[20*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:19*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[21*DATA_WIDTH-1:20*DATA_WIDTH] = valid_force_values[21*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:20*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[22*DATA_WIDTH-1:21*DATA_WIDTH] = valid_force_values[22*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:21*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[23*DATA_WIDTH-1:22*DATA_WIDTH] = valid_force_values[23*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:22*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[24*DATA_WIDTH-1:23*DATA_WIDTH] = valid_force_values[24*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:23*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[25*DATA_WIDTH-1:24*DATA_WIDTH] = valid_force_values[25*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:24*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[26*DATA_WIDTH-1:25*DATA_WIDTH] = valid_force_values[26*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:25*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[27*DATA_WIDTH-1:26*DATA_WIDTH] = valid_force_values[27*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:26*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[28*DATA_WIDTH-1:27*DATA_WIDTH] = valid_force_values[28*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:27*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[29*DATA_WIDTH-1:28*DATA_WIDTH] = valid_force_values[29*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:28*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[30*DATA_WIDTH-1:29*DATA_WIDTH] = valid_force_values[30*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:29*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[31*DATA_WIDTH-1:30*DATA_WIDTH] = valid_force_values[31*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:30*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[32*DATA_WIDTH-1:31*DATA_WIDTH] = valid_force_values[32*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:31*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[33*DATA_WIDTH-1:32*DATA_WIDTH] = valid_force_values[33*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:32*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[34*DATA_WIDTH-1:33*DATA_WIDTH] = valid_force_values[34*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:33*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[35*DATA_WIDTH-1:34*DATA_WIDTH] = valid_force_values[35*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:34*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[36*DATA_WIDTH-1:35*DATA_WIDTH] = valid_force_values[36*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:35*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[37*DATA_WIDTH-1:36*DATA_WIDTH] = valid_force_values[37*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:36*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[38*DATA_WIDTH-1:37*DATA_WIDTH] = valid_force_values[38*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:37*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[39*DATA_WIDTH-1:38*DATA_WIDTH] = valid_force_values[39*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:38*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[40*DATA_WIDTH-1:39*DATA_WIDTH] = valid_force_values[40*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:39*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[41*DATA_WIDTH-1:40*DATA_WIDTH] = valid_force_values[41*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:40*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[42*DATA_WIDTH-1:41*DATA_WIDTH] = valid_force_values[42*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:41*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[43*DATA_WIDTH-1:42*DATA_WIDTH] = valid_force_values[43*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:42*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[44*DATA_WIDTH-1:43*DATA_WIDTH] = valid_force_values[44*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:43*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[45*DATA_WIDTH-1:44*DATA_WIDTH] = valid_force_values[45*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:44*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[46*DATA_WIDTH-1:45*DATA_WIDTH] = valid_force_values[46*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:45*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[47*DATA_WIDTH-1:46*DATA_WIDTH] = valid_force_values[47*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:46*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[48*DATA_WIDTH-1:47*DATA_WIDTH] = valid_force_values[48*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:47*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[49*DATA_WIDTH-1:48*DATA_WIDTH] = valid_force_values[49*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:48*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[50*DATA_WIDTH-1:49*DATA_WIDTH] = valid_force_values[50*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:49*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[51*DATA_WIDTH-1:50*DATA_WIDTH] = valid_force_values[51*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:50*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[52*DATA_WIDTH-1:51*DATA_WIDTH] = valid_force_values[52*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:51*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[53*DATA_WIDTH-1:52*DATA_WIDTH] = valid_force_values[53*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:52*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[54*DATA_WIDTH-1:53*DATA_WIDTH] = valid_force_values[54*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:53*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[55*DATA_WIDTH-1:54*DATA_WIDTH] = valid_force_values[55*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:54*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[56*DATA_WIDTH-1:55*DATA_WIDTH] = valid_force_values[56*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:55*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[57*DATA_WIDTH-1:56*DATA_WIDTH] = valid_force_values[57*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:56*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[58*DATA_WIDTH-1:57*DATA_WIDTH] = valid_force_values[58*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:57*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[59*DATA_WIDTH-1:58*DATA_WIDTH] = valid_force_values[59*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:58*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[60*DATA_WIDTH-1:59*DATA_WIDTH] = valid_force_values[60*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:59*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[61*DATA_WIDTH-1:60*DATA_WIDTH] = valid_force_values[61*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:60*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[62*DATA_WIDTH-1:61*DATA_WIDTH] = valid_force_values[62*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:61*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[63*DATA_WIDTH-1:62*DATA_WIDTH] = valid_force_values[63*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:62*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	assign to_force_cache_LJ_Force_X[64*DATA_WIDTH-1:63*DATA_WIDTH] = valid_force_values[64*FORCE_EVAL_FIFO_DATA_WIDTH-2*DATA_WIDTH-1:63*FORCE_EVAL_FIFO_DATA_WIDTH+PARTICLE_ID_WIDTH+1];
	
	assign to_force_cache_particle_id[1*PARTICLE_ID_WIDTH-1:0*PARTICLE_ID_WIDTH] = valid_force_values[1*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:0*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[2*PARTICLE_ID_WIDTH-1:1*PARTICLE_ID_WIDTH] = valid_force_values[2*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:1*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[3*PARTICLE_ID_WIDTH-1:2*PARTICLE_ID_WIDTH] = valid_force_values[3*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:2*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[4*PARTICLE_ID_WIDTH-1:3*PARTICLE_ID_WIDTH] = valid_force_values[4*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:3*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[5*PARTICLE_ID_WIDTH-1:4*PARTICLE_ID_WIDTH] = valid_force_values[5*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:4*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[6*PARTICLE_ID_WIDTH-1:5*PARTICLE_ID_WIDTH] = valid_force_values[6*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:5*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[7*PARTICLE_ID_WIDTH-1:6*PARTICLE_ID_WIDTH] = valid_force_values[7*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:6*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[8*PARTICLE_ID_WIDTH-1:7*PARTICLE_ID_WIDTH] = valid_force_values[8*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:7*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[9*PARTICLE_ID_WIDTH-1:8*PARTICLE_ID_WIDTH] = valid_force_values[9*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:8*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[10*PARTICLE_ID_WIDTH-1:9*PARTICLE_ID_WIDTH] = valid_force_values[10*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:9*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[11*PARTICLE_ID_WIDTH-1:10*PARTICLE_ID_WIDTH] = valid_force_values[11*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:10*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[12*PARTICLE_ID_WIDTH-1:11*PARTICLE_ID_WIDTH] = valid_force_values[12*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:11*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[13*PARTICLE_ID_WIDTH-1:12*PARTICLE_ID_WIDTH] = valid_force_values[13*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:12*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[14*PARTICLE_ID_WIDTH-1:13*PARTICLE_ID_WIDTH] = valid_force_values[14*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:13*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[15*PARTICLE_ID_WIDTH-1:14*PARTICLE_ID_WIDTH] = valid_force_values[15*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:14*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[16*PARTICLE_ID_WIDTH-1:15*PARTICLE_ID_WIDTH] = valid_force_values[16*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:15*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[17*PARTICLE_ID_WIDTH-1:16*PARTICLE_ID_WIDTH] = valid_force_values[17*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:16*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[18*PARTICLE_ID_WIDTH-1:17*PARTICLE_ID_WIDTH] = valid_force_values[18*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:17*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[19*PARTICLE_ID_WIDTH-1:18*PARTICLE_ID_WIDTH] = valid_force_values[19*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:18*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[20*PARTICLE_ID_WIDTH-1:19*PARTICLE_ID_WIDTH] = valid_force_values[20*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:19*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[21*PARTICLE_ID_WIDTH-1:20*PARTICLE_ID_WIDTH] = valid_force_values[21*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:20*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[22*PARTICLE_ID_WIDTH-1:21*PARTICLE_ID_WIDTH] = valid_force_values[22*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:21*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[23*PARTICLE_ID_WIDTH-1:22*PARTICLE_ID_WIDTH] = valid_force_values[23*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:22*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[24*PARTICLE_ID_WIDTH-1:23*PARTICLE_ID_WIDTH] = valid_force_values[24*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:23*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[25*PARTICLE_ID_WIDTH-1:24*PARTICLE_ID_WIDTH] = valid_force_values[25*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:24*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[26*PARTICLE_ID_WIDTH-1:25*PARTICLE_ID_WIDTH] = valid_force_values[26*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:25*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[27*PARTICLE_ID_WIDTH-1:26*PARTICLE_ID_WIDTH] = valid_force_values[27*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:26*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[28*PARTICLE_ID_WIDTH-1:27*PARTICLE_ID_WIDTH] = valid_force_values[28*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:27*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[29*PARTICLE_ID_WIDTH-1:28*PARTICLE_ID_WIDTH] = valid_force_values[29*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:28*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[30*PARTICLE_ID_WIDTH-1:29*PARTICLE_ID_WIDTH] = valid_force_values[30*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:29*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[31*PARTICLE_ID_WIDTH-1:30*PARTICLE_ID_WIDTH] = valid_force_values[31*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:30*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[32*PARTICLE_ID_WIDTH-1:31*PARTICLE_ID_WIDTH] = valid_force_values[32*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:31*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[33*PARTICLE_ID_WIDTH-1:32*PARTICLE_ID_WIDTH] = valid_force_values[33*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:32*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[34*PARTICLE_ID_WIDTH-1:33*PARTICLE_ID_WIDTH] = valid_force_values[34*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:33*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[35*PARTICLE_ID_WIDTH-1:34*PARTICLE_ID_WIDTH] = valid_force_values[35*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:34*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[36*PARTICLE_ID_WIDTH-1:35*PARTICLE_ID_WIDTH] = valid_force_values[36*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:35*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[37*PARTICLE_ID_WIDTH-1:36*PARTICLE_ID_WIDTH] = valid_force_values[37*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:36*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[38*PARTICLE_ID_WIDTH-1:37*PARTICLE_ID_WIDTH] = valid_force_values[38*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:37*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[39*PARTICLE_ID_WIDTH-1:38*PARTICLE_ID_WIDTH] = valid_force_values[39*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:38*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[40*PARTICLE_ID_WIDTH-1:39*PARTICLE_ID_WIDTH] = valid_force_values[40*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:39*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[41*PARTICLE_ID_WIDTH-1:40*PARTICLE_ID_WIDTH] = valid_force_values[41*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:40*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[42*PARTICLE_ID_WIDTH-1:41*PARTICLE_ID_WIDTH] = valid_force_values[42*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:41*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[43*PARTICLE_ID_WIDTH-1:42*PARTICLE_ID_WIDTH] = valid_force_values[43*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:42*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[44*PARTICLE_ID_WIDTH-1:43*PARTICLE_ID_WIDTH] = valid_force_values[44*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:43*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[45*PARTICLE_ID_WIDTH-1:44*PARTICLE_ID_WIDTH] = valid_force_values[45*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:44*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[46*PARTICLE_ID_WIDTH-1:45*PARTICLE_ID_WIDTH] = valid_force_values[46*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:45*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[47*PARTICLE_ID_WIDTH-1:46*PARTICLE_ID_WIDTH] = valid_force_values[47*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:46*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[48*PARTICLE_ID_WIDTH-1:47*PARTICLE_ID_WIDTH] = valid_force_values[48*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:47*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[49*PARTICLE_ID_WIDTH-1:48*PARTICLE_ID_WIDTH] = valid_force_values[49*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:48*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[50*PARTICLE_ID_WIDTH-1:49*PARTICLE_ID_WIDTH] = valid_force_values[50*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:49*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[51*PARTICLE_ID_WIDTH-1:50*PARTICLE_ID_WIDTH] = valid_force_values[51*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:50*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[52*PARTICLE_ID_WIDTH-1:51*PARTICLE_ID_WIDTH] = valid_force_values[52*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:51*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[53*PARTICLE_ID_WIDTH-1:52*PARTICLE_ID_WIDTH] = valid_force_values[53*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:52*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[54*PARTICLE_ID_WIDTH-1:53*PARTICLE_ID_WIDTH] = valid_force_values[54*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:53*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[55*PARTICLE_ID_WIDTH-1:54*PARTICLE_ID_WIDTH] = valid_force_values[55*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:54*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[56*PARTICLE_ID_WIDTH-1:55*PARTICLE_ID_WIDTH] = valid_force_values[56*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:55*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[57*PARTICLE_ID_WIDTH-1:56*PARTICLE_ID_WIDTH] = valid_force_values[57*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:56*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[58*PARTICLE_ID_WIDTH-1:57*PARTICLE_ID_WIDTH] = valid_force_values[58*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:57*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[59*PARTICLE_ID_WIDTH-1:58*PARTICLE_ID_WIDTH] = valid_force_values[59*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:58*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[60*PARTICLE_ID_WIDTH-1:59*PARTICLE_ID_WIDTH] = valid_force_values[60*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:59*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[61*PARTICLE_ID_WIDTH-1:60*PARTICLE_ID_WIDTH] = valid_force_values[61*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:60*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[62*PARTICLE_ID_WIDTH-1:61*PARTICLE_ID_WIDTH] = valid_force_values[62*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:61*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[63*PARTICLE_ID_WIDTH-1:62*PARTICLE_ID_WIDTH] = valid_force_values[63*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:62*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	assign to_force_cache_particle_id[64*PARTICLE_ID_WIDTH-1:63*PARTICLE_ID_WIDTH] = valid_force_values[64*FORCE_EVAL_FIFO_DATA_WIDTH-3*DATA_WIDTH-1:63*FORCE_EVAL_FIFO_DATA_WIDTH+1];
	
	assign to_force_cache_partial_force_valid[0] = valid_force_values[0*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[1] = valid_force_values[1*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[2] = valid_force_values[2*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[3] = valid_force_values[3*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[4] = valid_force_values[4*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[5] = valid_force_values[5*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[6] = valid_force_values[6*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[7] = valid_force_values[7*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[8] = valid_force_values[8*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[9] = valid_force_values[9*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[10] = valid_force_values[10*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[11] = valid_force_values[11*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[12] = valid_force_values[12*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[13] = valid_force_values[13*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[14] = valid_force_values[14*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[15] = valid_force_values[15*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[16] = valid_force_values[16*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[17] = valid_force_values[17*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[18] = valid_force_values[18*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[19] = valid_force_values[19*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[20] = valid_force_values[20*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[21] = valid_force_values[21*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[22] = valid_force_values[22*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[23] = valid_force_values[23*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[24] = valid_force_values[24*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[25] = valid_force_values[25*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[26] = valid_force_values[26*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[27] = valid_force_values[27*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[28] = valid_force_values[28*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[29] = valid_force_values[29*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[30] = valid_force_values[30*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[31] = valid_force_values[31*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[32] = valid_force_values[32*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[33] = valid_force_values[33*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[34] = valid_force_values[34*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[35] = valid_force_values[35*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[36] = valid_force_values[36*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[37] = valid_force_values[37*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[38] = valid_force_values[38*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[39] = valid_force_values[39*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[40] = valid_force_values[40*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[41] = valid_force_values[41*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[42] = valid_force_values[42*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[43] = valid_force_values[43*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[44] = valid_force_values[44*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[45] = valid_force_values[45*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[46] = valid_force_values[46*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[47] = valid_force_values[47*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[48] = valid_force_values[48*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[49] = valid_force_values[49*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[50] = valid_force_values[50*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[51] = valid_force_values[51*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[52] = valid_force_values[52*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[53] = valid_force_values[53*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[54] = valid_force_values[54*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[55] = valid_force_values[55*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[56] = valid_force_values[56*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[57] = valid_force_values[57*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[58] = valid_force_values[58*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[59] = valid_force_values[59*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[60] = valid_force_values[60*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[61] = valid_force_values[61*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[62] = valid_force_values[62*FORCE_EVAL_FIFO_DATA_WIDTH];
	assign to_force_cache_partial_force_valid[63] = valid_force_values[63*FORCE_EVAL_FIFO_DATA_WIDTH];
	// Force_Cache_1_1_1
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_1_1_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[0]),
		.in_particle_id(to_force_cache_particle_id[1*PARTICLE_ID_WIDTH-1:0*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[1*DATA_WIDTH-1:0*DATA_WIDTH], to_force_cache_LJ_Force_Y[1*DATA_WIDTH-1:0*DATA_WIDTH], to_force_cache_LJ_Force_X[1*DATA_WIDTH-1:0*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[0]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[1*PARTICLE_ID_WIDTH-1:0*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[0])
	);
	// Force_Cache_1_1_2
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_1_1_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[1]),
		.in_particle_id(to_force_cache_particle_id[2*PARTICLE_ID_WIDTH-1:1*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[2*DATA_WIDTH-1:1*DATA_WIDTH], to_force_cache_LJ_Force_Y[2*DATA_WIDTH-1:1*DATA_WIDTH], to_force_cache_LJ_Force_X[2*DATA_WIDTH-1:1*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[1]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[2*PARTICLE_ID_WIDTH-1:1*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[1])
	);
	// Force_Cache_1_1_3
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_1_1_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[2]),
		.in_particle_id(to_force_cache_particle_id[3*PARTICLE_ID_WIDTH-1:2*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[3*DATA_WIDTH-1:2*DATA_WIDTH], to_force_cache_LJ_Force_Y[3*DATA_WIDTH-1:2*DATA_WIDTH], to_force_cache_LJ_Force_X[3*DATA_WIDTH-1:2*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[2]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[3*PARTICLE_ID_WIDTH-1:2*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[2])
	);
	// Force_Cache_1_1_4
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_1_1_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[3]),
		.in_particle_id(to_force_cache_particle_id[4*PARTICLE_ID_WIDTH-1:3*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[4*DATA_WIDTH-1:3*DATA_WIDTH], to_force_cache_LJ_Force_Y[4*DATA_WIDTH-1:3*DATA_WIDTH], to_force_cache_LJ_Force_X[4*DATA_WIDTH-1:3*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[3]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[4*PARTICLE_ID_WIDTH-1:3*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[3])
	);
	// Force_Cache_1_2_1
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_1_2_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[4]),
		.in_particle_id(to_force_cache_particle_id[5*PARTICLE_ID_WIDTH-1:4*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[5*DATA_WIDTH-1:4*DATA_WIDTH], to_force_cache_LJ_Force_Y[5*DATA_WIDTH-1:4*DATA_WIDTH], to_force_cache_LJ_Force_X[5*DATA_WIDTH-1:4*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[4]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[5*PARTICLE_ID_WIDTH-1:4*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[4])
	);
	// Force_Cache_1_2_2
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_1_2_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[5]),
		.in_particle_id(to_force_cache_particle_id[6*PARTICLE_ID_WIDTH-1:5*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[6*DATA_WIDTH-1:5*DATA_WIDTH], to_force_cache_LJ_Force_Y[6*DATA_WIDTH-1:5*DATA_WIDTH], to_force_cache_LJ_Force_X[6*DATA_WIDTH-1:5*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[5]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[6*PARTICLE_ID_WIDTH-1:5*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[5])
	);
	// Force_Cache_1_2_3
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_1_2_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[6]),
		.in_particle_id(to_force_cache_particle_id[7*PARTICLE_ID_WIDTH-1:6*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[7*DATA_WIDTH-1:6*DATA_WIDTH], to_force_cache_LJ_Force_Y[7*DATA_WIDTH-1:6*DATA_WIDTH], to_force_cache_LJ_Force_X[7*DATA_WIDTH-1:6*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[6]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[7*PARTICLE_ID_WIDTH-1:6*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[6])
	);
	// Force_Cache_1_2_4
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_1_2_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[7]),
		.in_particle_id(to_force_cache_particle_id[8*PARTICLE_ID_WIDTH-1:7*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[8*DATA_WIDTH-1:7*DATA_WIDTH], to_force_cache_LJ_Force_Y[8*DATA_WIDTH-1:7*DATA_WIDTH], to_force_cache_LJ_Force_X[8*DATA_WIDTH-1:7*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[7]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[8*PARTICLE_ID_WIDTH-1:7*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[7])
	);
	// Force_Cache_1_3_1
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_1_3_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[8]),
		.in_particle_id(to_force_cache_particle_id[9*PARTICLE_ID_WIDTH-1:8*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[9*DATA_WIDTH-1:8*DATA_WIDTH], to_force_cache_LJ_Force_Y[9*DATA_WIDTH-1:8*DATA_WIDTH], to_force_cache_LJ_Force_X[9*DATA_WIDTH-1:8*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[8]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[9*3*DATA_WIDTH-1:8*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[9*PARTICLE_ID_WIDTH-1:8*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[8])
	);
	// Force_Cache_1_3_2
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_1_3_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[9]),
		.in_particle_id(to_force_cache_particle_id[10*PARTICLE_ID_WIDTH-1:9*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[10*DATA_WIDTH-1:9*DATA_WIDTH], to_force_cache_LJ_Force_Y[10*DATA_WIDTH-1:9*DATA_WIDTH], to_force_cache_LJ_Force_X[10*DATA_WIDTH-1:9*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[9]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[10*3*DATA_WIDTH-1:9*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[10*PARTICLE_ID_WIDTH-1:9*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[9])
	);
	// Force_Cache_1_3_3
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_1_3_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[10]),
		.in_particle_id(to_force_cache_particle_id[11*PARTICLE_ID_WIDTH-1:10*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[11*DATA_WIDTH-1:10*DATA_WIDTH], to_force_cache_LJ_Force_Y[11*DATA_WIDTH-1:10*DATA_WIDTH], to_force_cache_LJ_Force_X[11*DATA_WIDTH-1:10*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[10]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[11*3*DATA_WIDTH-1:10*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[11*PARTICLE_ID_WIDTH-1:10*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[10])
	);
	// Force_Cache_1_3_4
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_1_3_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[11]),
		.in_particle_id(to_force_cache_particle_id[12*PARTICLE_ID_WIDTH-1:11*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[12*DATA_WIDTH-1:11*DATA_WIDTH], to_force_cache_LJ_Force_Y[12*DATA_WIDTH-1:11*DATA_WIDTH], to_force_cache_LJ_Force_X[12*DATA_WIDTH-1:11*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[11]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[12*3*DATA_WIDTH-1:11*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[12*PARTICLE_ID_WIDTH-1:11*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[11])
	);
	// Force_Cache_1_4_1
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_1_4_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[12]),
		.in_particle_id(to_force_cache_particle_id[13*PARTICLE_ID_WIDTH-1:12*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[13*DATA_WIDTH-1:12*DATA_WIDTH], to_force_cache_LJ_Force_Y[13*DATA_WIDTH-1:12*DATA_WIDTH], to_force_cache_LJ_Force_X[13*DATA_WIDTH-1:12*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[12]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[13*3*DATA_WIDTH-1:12*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[13*PARTICLE_ID_WIDTH-1:12*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[12])
	);
	// Force_Cache_1_4_2
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_1_4_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[13]),
		.in_particle_id(to_force_cache_particle_id[14*PARTICLE_ID_WIDTH-1:13*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[14*DATA_WIDTH-1:13*DATA_WIDTH], to_force_cache_LJ_Force_Y[14*DATA_WIDTH-1:13*DATA_WIDTH], to_force_cache_LJ_Force_X[14*DATA_WIDTH-1:13*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[13]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[14*3*DATA_WIDTH-1:13*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[14*PARTICLE_ID_WIDTH-1:13*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[13])
	);
	// Force_Cache_1_4_3
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_1_4_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[14]),
		.in_particle_id(to_force_cache_particle_id[15*PARTICLE_ID_WIDTH-1:14*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[15*DATA_WIDTH-1:14*DATA_WIDTH], to_force_cache_LJ_Force_Y[15*DATA_WIDTH-1:14*DATA_WIDTH], to_force_cache_LJ_Force_X[15*DATA_WIDTH-1:14*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[14]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[15*3*DATA_WIDTH-1:14*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[15*PARTICLE_ID_WIDTH-1:14*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[14])
	);
	// Force_Cache_1_4_4
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_1_4_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[15]),
		.in_particle_id(to_force_cache_particle_id[16*PARTICLE_ID_WIDTH-1:15*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[16*DATA_WIDTH-1:15*DATA_WIDTH], to_force_cache_LJ_Force_Y[16*DATA_WIDTH-1:15*DATA_WIDTH], to_force_cache_LJ_Force_X[16*DATA_WIDTH-1:15*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[15]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[16*3*DATA_WIDTH-1:15*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[16*PARTICLE_ID_WIDTH-1:15*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[15])
	);
	// Force_Cache_2_1_1
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_2_1_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[16]),
		.in_particle_id(to_force_cache_particle_id[17*PARTICLE_ID_WIDTH-1:16*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[17*DATA_WIDTH-1:16*DATA_WIDTH], to_force_cache_LJ_Force_Y[17*DATA_WIDTH-1:16*DATA_WIDTH], to_force_cache_LJ_Force_X[17*DATA_WIDTH-1:16*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[16]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[17*PARTICLE_ID_WIDTH-1:16*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[16])
	);
	// Force_Cache_2_1_2
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_2_1_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[17]),
		.in_particle_id(to_force_cache_particle_id[18*PARTICLE_ID_WIDTH-1:17*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[18*DATA_WIDTH-1:17*DATA_WIDTH], to_force_cache_LJ_Force_Y[18*DATA_WIDTH-1:17*DATA_WIDTH], to_force_cache_LJ_Force_X[18*DATA_WIDTH-1:17*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[17]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[18*PARTICLE_ID_WIDTH-1:17*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[17])
	);
	// Force_Cache_2_1_3
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_2_1_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[18]),
		.in_particle_id(to_force_cache_particle_id[19*PARTICLE_ID_WIDTH-1:18*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[19*DATA_WIDTH-1:18*DATA_WIDTH], to_force_cache_LJ_Force_Y[19*DATA_WIDTH-1:18*DATA_WIDTH], to_force_cache_LJ_Force_X[19*DATA_WIDTH-1:18*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[18]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[19*PARTICLE_ID_WIDTH-1:18*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[18])
	);
	// Force_Cache_2_1_4
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_2_1_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[19]),
		.in_particle_id(to_force_cache_particle_id[20*PARTICLE_ID_WIDTH-1:19*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[20*DATA_WIDTH-1:19*DATA_WIDTH], to_force_cache_LJ_Force_Y[20*DATA_WIDTH-1:19*DATA_WIDTH], to_force_cache_LJ_Force_X[20*DATA_WIDTH-1:19*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[19]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[20*PARTICLE_ID_WIDTH-1:19*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[19])
	);
	// Force_Cache_2_2_1
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_2_2_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[20]),
		.in_particle_id(to_force_cache_particle_id[21*PARTICLE_ID_WIDTH-1:20*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[21*DATA_WIDTH-1:20*DATA_WIDTH], to_force_cache_LJ_Force_Y[21*DATA_WIDTH-1:20*DATA_WIDTH], to_force_cache_LJ_Force_X[21*DATA_WIDTH-1:20*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[20]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[21*PARTICLE_ID_WIDTH-1:20*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[20])
	);
	// Force_Cache_2_2_2
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_2_2_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[21]),
		.in_particle_id(to_force_cache_particle_id[22*PARTICLE_ID_WIDTH-1:21*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[22*DATA_WIDTH-1:21*DATA_WIDTH], to_force_cache_LJ_Force_Y[22*DATA_WIDTH-1:21*DATA_WIDTH], to_force_cache_LJ_Force_X[22*DATA_WIDTH-1:21*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[21]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[22*PARTICLE_ID_WIDTH-1:21*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[21])
	);
	// Force_Cache_2_2_3
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_2_2_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[22]),
		.in_particle_id(to_force_cache_particle_id[23*PARTICLE_ID_WIDTH-1:22*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[23*DATA_WIDTH-1:22*DATA_WIDTH], to_force_cache_LJ_Force_Y[23*DATA_WIDTH-1:22*DATA_WIDTH], to_force_cache_LJ_Force_X[23*DATA_WIDTH-1:22*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[22]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[23*PARTICLE_ID_WIDTH-1:22*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[22])
	);
	// Force_Cache_2_2_4
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_2_2_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[23]),
		.in_particle_id(to_force_cache_particle_id[24*PARTICLE_ID_WIDTH-1:23*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[24*DATA_WIDTH-1:23*DATA_WIDTH], to_force_cache_LJ_Force_Y[24*DATA_WIDTH-1:23*DATA_WIDTH], to_force_cache_LJ_Force_X[24*DATA_WIDTH-1:23*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[23]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[24*PARTICLE_ID_WIDTH-1:23*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[23])
	);
	// Force_Cache_2_3_1
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_2_3_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[24]),
		.in_particle_id(to_force_cache_particle_id[25*PARTICLE_ID_WIDTH-1:24*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[25*DATA_WIDTH-1:24*DATA_WIDTH], to_force_cache_LJ_Force_Y[25*DATA_WIDTH-1:24*DATA_WIDTH], to_force_cache_LJ_Force_X[25*DATA_WIDTH-1:24*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[24]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[25*3*DATA_WIDTH-1:24*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[25*PARTICLE_ID_WIDTH-1:24*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[24])
	);
	// Force_Cache_2_3_2
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_2_3_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[25]),
		.in_particle_id(to_force_cache_particle_id[26*PARTICLE_ID_WIDTH-1:25*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[26*DATA_WIDTH-1:25*DATA_WIDTH], to_force_cache_LJ_Force_Y[26*DATA_WIDTH-1:25*DATA_WIDTH], to_force_cache_LJ_Force_X[26*DATA_WIDTH-1:25*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[25]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[26*3*DATA_WIDTH-1:25*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[26*PARTICLE_ID_WIDTH-1:25*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[25])
	);
	// Force_Cache_2_3_3
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_2_3_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[26]),
		.in_particle_id(to_force_cache_particle_id[27*PARTICLE_ID_WIDTH-1:26*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[27*DATA_WIDTH-1:26*DATA_WIDTH], to_force_cache_LJ_Force_Y[27*DATA_WIDTH-1:26*DATA_WIDTH], to_force_cache_LJ_Force_X[27*DATA_WIDTH-1:26*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[26]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[27*3*DATA_WIDTH-1:26*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[27*PARTICLE_ID_WIDTH-1:26*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[26])
	);
	// Force_Cache_2_3_4
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_2_3_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[27]),
		.in_particle_id(to_force_cache_particle_id[28*PARTICLE_ID_WIDTH-1:27*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[28*DATA_WIDTH-1:27*DATA_WIDTH], to_force_cache_LJ_Force_Y[28*DATA_WIDTH-1:27*DATA_WIDTH], to_force_cache_LJ_Force_X[28*DATA_WIDTH-1:27*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[27]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[28*3*DATA_WIDTH-1:27*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[28*PARTICLE_ID_WIDTH-1:27*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[27])
	);
	// Force_Cache_2_4_1
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_2_4_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[28]),
		.in_particle_id(to_force_cache_particle_id[29*PARTICLE_ID_WIDTH-1:28*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[29*DATA_WIDTH-1:28*DATA_WIDTH], to_force_cache_LJ_Force_Y[29*DATA_WIDTH-1:28*DATA_WIDTH], to_force_cache_LJ_Force_X[29*DATA_WIDTH-1:28*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[28]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[29*PARTICLE_ID_WIDTH-1:28*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[28])
	);
	// Force_Cache_2_4_2
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_2_4_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[29]),
		.in_particle_id(to_force_cache_particle_id[30*PARTICLE_ID_WIDTH-1:29*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[30*DATA_WIDTH-1:29*DATA_WIDTH], to_force_cache_LJ_Force_Y[30*DATA_WIDTH-1:29*DATA_WIDTH], to_force_cache_LJ_Force_X[30*DATA_WIDTH-1:29*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[29]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[30*PARTICLE_ID_WIDTH-1:29*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[29])
	);
	// Force_Cache_2_4_3
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_2_4_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[30]),
		.in_particle_id(to_force_cache_particle_id[31*PARTICLE_ID_WIDTH-1:30*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[31*DATA_WIDTH-1:30*DATA_WIDTH], to_force_cache_LJ_Force_Y[31*DATA_WIDTH-1:30*DATA_WIDTH], to_force_cache_LJ_Force_X[31*DATA_WIDTH-1:30*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[30]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[31*PARTICLE_ID_WIDTH-1:30*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[30])
	);
	// Force_Cache_2_4_4
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_2_4_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[31]),
		.in_particle_id(to_force_cache_particle_id[32*PARTICLE_ID_WIDTH-1:31*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[32*DATA_WIDTH-1:31*DATA_WIDTH], to_force_cache_LJ_Force_Y[32*DATA_WIDTH-1:31*DATA_WIDTH], to_force_cache_LJ_Force_X[32*DATA_WIDTH-1:31*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[31]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[32*PARTICLE_ID_WIDTH-1:31*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[31])
	);
	// Force_Cache_3_1_1
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_3_1_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[32]),
		.in_particle_id(to_force_cache_particle_id[33*PARTICLE_ID_WIDTH-1:32*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[33*DATA_WIDTH-1:32*DATA_WIDTH], to_force_cache_LJ_Force_Y[33*DATA_WIDTH-1:32*DATA_WIDTH], to_force_cache_LJ_Force_X[33*DATA_WIDTH-1:32*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[32]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[33*3*DATA_WIDTH-1:32*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[33*PARTICLE_ID_WIDTH-1:32*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[32])
	);
	// Force_Cache_3_1_2
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_3_1_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[33]),
		.in_particle_id(to_force_cache_particle_id[34*PARTICLE_ID_WIDTH-1:33*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[34*DATA_WIDTH-1:33*DATA_WIDTH], to_force_cache_LJ_Force_Y[34*DATA_WIDTH-1:33*DATA_WIDTH], to_force_cache_LJ_Force_X[34*DATA_WIDTH-1:33*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[33]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[34*3*DATA_WIDTH-1:33*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[34*PARTICLE_ID_WIDTH-1:33*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[33])
	);
	// Force_Cache_3_1_3
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_3_1_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[34]),
		.in_particle_id(to_force_cache_particle_id[35*PARTICLE_ID_WIDTH-1:34*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[35*DATA_WIDTH-1:34*DATA_WIDTH], to_force_cache_LJ_Force_Y[35*DATA_WIDTH-1:34*DATA_WIDTH], to_force_cache_LJ_Force_X[35*DATA_WIDTH-1:34*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[34]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[35*3*DATA_WIDTH-1:34*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[35*PARTICLE_ID_WIDTH-1:34*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[34])
	);
	// Force_Cache_3_1_4
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_3_1_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[35]),
		.in_particle_id(to_force_cache_particle_id[36*PARTICLE_ID_WIDTH-1:35*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[36*DATA_WIDTH-1:35*DATA_WIDTH], to_force_cache_LJ_Force_Y[36*DATA_WIDTH-1:35*DATA_WIDTH], to_force_cache_LJ_Force_X[36*DATA_WIDTH-1:35*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[35]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[36*3*DATA_WIDTH-1:35*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[36*PARTICLE_ID_WIDTH-1:35*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[35])
	);
	// Force_Cache_3_2_1
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_3_2_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[36]),
		.in_particle_id(to_force_cache_particle_id[37*PARTICLE_ID_WIDTH-1:36*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[37*DATA_WIDTH-1:36*DATA_WIDTH], to_force_cache_LJ_Force_Y[37*DATA_WIDTH-1:36*DATA_WIDTH], to_force_cache_LJ_Force_X[37*DATA_WIDTH-1:36*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[36]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[37*3*DATA_WIDTH-1:36*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[37*PARTICLE_ID_WIDTH-1:36*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[36])
	);
	// Force_Cache_3_2_2
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_3_2_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[37]),
		.in_particle_id(to_force_cache_particle_id[38*PARTICLE_ID_WIDTH-1:37*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[38*DATA_WIDTH-1:37*DATA_WIDTH], to_force_cache_LJ_Force_Y[38*DATA_WIDTH-1:37*DATA_WIDTH], to_force_cache_LJ_Force_X[38*DATA_WIDTH-1:37*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[37]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[38*3*DATA_WIDTH-1:37*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[38*PARTICLE_ID_WIDTH-1:37*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[37])
	);
	// Force_Cache_3_2_3
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_3_2_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[38]),
		.in_particle_id(to_force_cache_particle_id[39*PARTICLE_ID_WIDTH-1:38*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[39*DATA_WIDTH-1:38*DATA_WIDTH], to_force_cache_LJ_Force_Y[39*DATA_WIDTH-1:38*DATA_WIDTH], to_force_cache_LJ_Force_X[39*DATA_WIDTH-1:38*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[38]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[39*3*DATA_WIDTH-1:38*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[39*PARTICLE_ID_WIDTH-1:38*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[38])
	);
	// Force_Cache_3_2_4
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_3_2_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[39]),
		.in_particle_id(to_force_cache_particle_id[40*PARTICLE_ID_WIDTH-1:39*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[40*DATA_WIDTH-1:39*DATA_WIDTH], to_force_cache_LJ_Force_Y[40*DATA_WIDTH-1:39*DATA_WIDTH], to_force_cache_LJ_Force_X[40*DATA_WIDTH-1:39*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[39]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[40*3*DATA_WIDTH-1:39*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[40*PARTICLE_ID_WIDTH-1:39*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[39])
	);
	// Force_Cache_3_3_1
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_3_3_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[40]),
		.in_particle_id(to_force_cache_particle_id[41*PARTICLE_ID_WIDTH-1:40*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[41*DATA_WIDTH-1:40*DATA_WIDTH], to_force_cache_LJ_Force_Y[41*DATA_WIDTH-1:40*DATA_WIDTH], to_force_cache_LJ_Force_X[41*DATA_WIDTH-1:40*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[40]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[41*3*DATA_WIDTH-1:40*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[41*PARTICLE_ID_WIDTH-1:40*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[40])
	);
	// Force_Cache_3_3_2
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_3_3_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[41]),
		.in_particle_id(to_force_cache_particle_id[42*PARTICLE_ID_WIDTH-1:41*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[42*DATA_WIDTH-1:41*DATA_WIDTH], to_force_cache_LJ_Force_Y[42*DATA_WIDTH-1:41*DATA_WIDTH], to_force_cache_LJ_Force_X[42*DATA_WIDTH-1:41*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[41]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[42*3*DATA_WIDTH-1:41*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[42*PARTICLE_ID_WIDTH-1:41*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[41])
	);
	// Force_Cache_3_3_3
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_3_3_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[42]),
		.in_particle_id(to_force_cache_particle_id[43*PARTICLE_ID_WIDTH-1:42*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[43*DATA_WIDTH-1:42*DATA_WIDTH], to_force_cache_LJ_Force_Y[43*DATA_WIDTH-1:42*DATA_WIDTH], to_force_cache_LJ_Force_X[43*DATA_WIDTH-1:42*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[42]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[43*3*DATA_WIDTH-1:42*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[43*PARTICLE_ID_WIDTH-1:42*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[42])
	);
	// Force_Cache_3_3_4
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_3_3_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[43]),
		.in_particle_id(to_force_cache_particle_id[44*PARTICLE_ID_WIDTH-1:43*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[44*DATA_WIDTH-1:43*DATA_WIDTH], to_force_cache_LJ_Force_Y[44*DATA_WIDTH-1:43*DATA_WIDTH], to_force_cache_LJ_Force_X[44*DATA_WIDTH-1:43*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[43]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[44*3*DATA_WIDTH-1:43*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[44*PARTICLE_ID_WIDTH-1:43*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[43])
	);
	// Force_Cache_3_4_1
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_3_4_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[44]),
		.in_particle_id(to_force_cache_particle_id[45*PARTICLE_ID_WIDTH-1:44*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[45*DATA_WIDTH-1:44*DATA_WIDTH], to_force_cache_LJ_Force_Y[45*DATA_WIDTH-1:44*DATA_WIDTH], to_force_cache_LJ_Force_X[45*DATA_WIDTH-1:44*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[44]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[45*3*DATA_WIDTH-1:44*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[45*PARTICLE_ID_WIDTH-1:44*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[44])
	);
	// Force_Cache_3_4_2
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_3_4_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[45]),
		.in_particle_id(to_force_cache_particle_id[46*PARTICLE_ID_WIDTH-1:45*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[46*DATA_WIDTH-1:45*DATA_WIDTH], to_force_cache_LJ_Force_Y[46*DATA_WIDTH-1:45*DATA_WIDTH], to_force_cache_LJ_Force_X[46*DATA_WIDTH-1:45*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[45]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[46*3*DATA_WIDTH-1:45*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[46*PARTICLE_ID_WIDTH-1:45*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[45])
	);
	// Force_Cache_3_4_3
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_3_4_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[46]),
		.in_particle_id(to_force_cache_particle_id[47*PARTICLE_ID_WIDTH-1:46*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[47*DATA_WIDTH-1:46*DATA_WIDTH], to_force_cache_LJ_Force_Y[47*DATA_WIDTH-1:46*DATA_WIDTH], to_force_cache_LJ_Force_X[47*DATA_WIDTH-1:46*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[46]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[47*3*DATA_WIDTH-1:46*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[47*PARTICLE_ID_WIDTH-1:46*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[46])
	);
	// Force_Cache_3_4_4
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_3_4_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[47]),
		.in_particle_id(to_force_cache_particle_id[48*PARTICLE_ID_WIDTH-1:47*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[48*DATA_WIDTH-1:47*DATA_WIDTH], to_force_cache_LJ_Force_Y[48*DATA_WIDTH-1:47*DATA_WIDTH], to_force_cache_LJ_Force_X[48*DATA_WIDTH-1:47*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[47]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[48*3*DATA_WIDTH-1:47*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[48*PARTICLE_ID_WIDTH-1:47*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[47])
	);
	// Force_Cache_4_1_1
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_4_1_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[48]),
		.in_particle_id(to_force_cache_particle_id[49*PARTICLE_ID_WIDTH-1:48*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[49*DATA_WIDTH-1:48*DATA_WIDTH], to_force_cache_LJ_Force_Y[49*DATA_WIDTH-1:48*DATA_WIDTH], to_force_cache_LJ_Force_X[49*DATA_WIDTH-1:48*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[48]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[49*3*DATA_WIDTH-1:48*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[49*PARTICLE_ID_WIDTH-1:48*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[48])
	);
	// Force_Cache_4_1_2
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_4_1_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[49]),
		.in_particle_id(to_force_cache_particle_id[50*PARTICLE_ID_WIDTH-1:49*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[50*DATA_WIDTH-1:49*DATA_WIDTH], to_force_cache_LJ_Force_Y[50*DATA_WIDTH-1:49*DATA_WIDTH], to_force_cache_LJ_Force_X[50*DATA_WIDTH-1:49*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[49]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[50*3*DATA_WIDTH-1:49*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[50*PARTICLE_ID_WIDTH-1:49*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[49])
	);
	// Force_Cache_4_1_3
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_4_1_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[50]),
		.in_particle_id(to_force_cache_particle_id[51*PARTICLE_ID_WIDTH-1:50*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[51*DATA_WIDTH-1:50*DATA_WIDTH], to_force_cache_LJ_Force_Y[51*DATA_WIDTH-1:50*DATA_WIDTH], to_force_cache_LJ_Force_X[51*DATA_WIDTH-1:50*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[50]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[51*3*DATA_WIDTH-1:50*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[51*PARTICLE_ID_WIDTH-1:50*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[50])
	);
	// Force_Cache_4_1_4
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_4_1_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[51]),
		.in_particle_id(to_force_cache_particle_id[52*PARTICLE_ID_WIDTH-1:51*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[52*DATA_WIDTH-1:51*DATA_WIDTH], to_force_cache_LJ_Force_Y[52*DATA_WIDTH-1:51*DATA_WIDTH], to_force_cache_LJ_Force_X[52*DATA_WIDTH-1:51*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[51]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[52*3*DATA_WIDTH-1:51*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[52*PARTICLE_ID_WIDTH-1:51*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[51])
	);
	// Force_Cache_4_2_1
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_4_2_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[52]),
		.in_particle_id(to_force_cache_particle_id[53*PARTICLE_ID_WIDTH-1:52*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[53*DATA_WIDTH-1:52*DATA_WIDTH], to_force_cache_LJ_Force_Y[53*DATA_WIDTH-1:52*DATA_WIDTH], to_force_cache_LJ_Force_X[53*DATA_WIDTH-1:52*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[52]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[53*3*DATA_WIDTH-1:52*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[53*PARTICLE_ID_WIDTH-1:52*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[52])
	);
	// Force_Cache_4_2_2
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_4_2_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[53]),
		.in_particle_id(to_force_cache_particle_id[54*PARTICLE_ID_WIDTH-1:53*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[54*DATA_WIDTH-1:53*DATA_WIDTH], to_force_cache_LJ_Force_Y[54*DATA_WIDTH-1:53*DATA_WIDTH], to_force_cache_LJ_Force_X[54*DATA_WIDTH-1:53*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[53]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[54*3*DATA_WIDTH-1:53*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[54*PARTICLE_ID_WIDTH-1:53*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[53])
	);
	// Force_Cache_4_2_3
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_4_2_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[54]),
		.in_particle_id(to_force_cache_particle_id[55*PARTICLE_ID_WIDTH-1:54*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[55*DATA_WIDTH-1:54*DATA_WIDTH], to_force_cache_LJ_Force_Y[55*DATA_WIDTH-1:54*DATA_WIDTH], to_force_cache_LJ_Force_X[55*DATA_WIDTH-1:54*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[54]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[55*3*DATA_WIDTH-1:54*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[55*PARTICLE_ID_WIDTH-1:54*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[54])
	);
	// Force_Cache_4_2_4
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_4_2_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[55]),
		.in_particle_id(to_force_cache_particle_id[56*PARTICLE_ID_WIDTH-1:55*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[56*DATA_WIDTH-1:55*DATA_WIDTH], to_force_cache_LJ_Force_Y[56*DATA_WIDTH-1:55*DATA_WIDTH], to_force_cache_LJ_Force_X[56*DATA_WIDTH-1:55*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[55]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[56*3*DATA_WIDTH-1:55*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[56*PARTICLE_ID_WIDTH-1:55*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[55])
	);
	// Force_Cache_4_3_1
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_4_3_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[56]),
		.in_particle_id(to_force_cache_particle_id[57*PARTICLE_ID_WIDTH-1:56*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[57*DATA_WIDTH-1:56*DATA_WIDTH], to_force_cache_LJ_Force_Y[57*DATA_WIDTH-1:56*DATA_WIDTH], to_force_cache_LJ_Force_X[57*DATA_WIDTH-1:56*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[56]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[57*3*DATA_WIDTH-1:56*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[57*PARTICLE_ID_WIDTH-1:56*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[56])
	);
	// Force_Cache_4_3_2
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_4_3_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[57]),
		.in_particle_id(to_force_cache_particle_id[58*PARTICLE_ID_WIDTH-1:57*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[58*DATA_WIDTH-1:57*DATA_WIDTH], to_force_cache_LJ_Force_Y[58*DATA_WIDTH-1:57*DATA_WIDTH], to_force_cache_LJ_Force_X[58*DATA_WIDTH-1:57*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[57]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[58*3*DATA_WIDTH-1:57*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[58*PARTICLE_ID_WIDTH-1:57*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[57])
	);
	// Force_Cache_4_3_3
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_4_3_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[58]),
		.in_particle_id(to_force_cache_particle_id[59*PARTICLE_ID_WIDTH-1:58*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[59*DATA_WIDTH-1:58*DATA_WIDTH], to_force_cache_LJ_Force_Y[59*DATA_WIDTH-1:58*DATA_WIDTH], to_force_cache_LJ_Force_X[59*DATA_WIDTH-1:58*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[58]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[59*3*DATA_WIDTH-1:58*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[59*PARTICLE_ID_WIDTH-1:58*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[58])
	);
	// Force_Cache_4_3_4
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_4_3_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[59]),
		.in_particle_id(to_force_cache_particle_id[60*PARTICLE_ID_WIDTH-1:59*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[60*DATA_WIDTH-1:59*DATA_WIDTH], to_force_cache_LJ_Force_Y[60*DATA_WIDTH-1:59*DATA_WIDTH], to_force_cache_LJ_Force_X[60*DATA_WIDTH-1:59*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[59]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[60*3*DATA_WIDTH-1:59*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[60*PARTICLE_ID_WIDTH-1:59*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[59])
	);
	// Force_Cache_4_4_1
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_4_4_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[60]),
		.in_particle_id(to_force_cache_particle_id[61*PARTICLE_ID_WIDTH-1:60*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[61*DATA_WIDTH-1:60*DATA_WIDTH], to_force_cache_LJ_Force_Y[61*DATA_WIDTH-1:60*DATA_WIDTH], to_force_cache_LJ_Force_X[61*DATA_WIDTH-1:60*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[60]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[61*3*DATA_WIDTH-1:60*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[61*PARTICLE_ID_WIDTH-1:60*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[60])
	);
	// Force_Cache_4_4_2
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_4_4_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[61]),
		.in_particle_id(to_force_cache_particle_id[62*PARTICLE_ID_WIDTH-1:61*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[62*DATA_WIDTH-1:61*DATA_WIDTH], to_force_cache_LJ_Force_Y[62*DATA_WIDTH-1:61*DATA_WIDTH], to_force_cache_LJ_Force_X[62*DATA_WIDTH-1:61*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[61]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[62*3*DATA_WIDTH-1:61*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[62*PARTICLE_ID_WIDTH-1:61*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[61])
	);
	// Force_Cache_4_4_3
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_4_4_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[62]),
		.in_particle_id(to_force_cache_particle_id[63*PARTICLE_ID_WIDTH-1:62*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[63*DATA_WIDTH-1:62*DATA_WIDTH], to_force_cache_LJ_Force_Y[63*DATA_WIDTH-1:62*DATA_WIDTH], to_force_cache_LJ_Force_X[63*DATA_WIDTH-1:62*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[62]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[63*3*DATA_WIDTH-1:62*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[63*PARTICLE_ID_WIDTH-1:62*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[62])
	);
	// Force_Cache_4_4_4
	Force_Write_Back_Controller_64_Cells
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Force_4_4_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(to_force_cache_partial_force_valid[63]),
		.in_particle_id(to_force_cache_particle_id[64*PARTICLE_ID_WIDTH-1:63*PARTICLE_ID_WIDTH]),
		.in_partial_force({to_force_cache_LJ_Force_Z[64*DATA_WIDTH-1:63*DATA_WIDTH], to_force_cache_LJ_Force_Y[64*DATA_WIDTH-1:63*DATA_WIDTH], to_force_cache_LJ_Force_X[64*DATA_WIDTH-1:63*DATA_WIDTH]}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[63]),									// Enables read data from the force cache, if this signal is high, then no write operation is permitted
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[64*3*DATA_WIDTH-1:63*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[64*PARTICLE_ID_WIDTH-1:63*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[63])
	);
	
endmodule