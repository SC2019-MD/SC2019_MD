/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Module: RL_LJ_Intergrated_Top.v
//
//	Function:
//				Integrated top module holding all the cells in the simulation space
//
//	Purpose:
//				For real simulation with all the dataset
//				Timing testing with the integrated system
//
// Data Organization:
//				Address 0 for each cell module: # of particles in the cell.
//				MSB-LSB: {posz, posy, posx}
//
// Used by:
//				NA
//
// Dependency:
//				RL_LJ_Evaluation_Unit.v
//				Particle_Pair_Gen_HalfShell.v
//				Motion_Update.v
//				cell_x_y_z.v
//				Force_Cache_x_y_z.v
//				Velocity_Cache_x_y_z.v
//
// Testbench:
//				TBD
//
// Timing:

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module RL_LJ_Intergrated_Top
#(
	parameter DATA_WIDTH 					= 32,
	// Simulation parameters
	parameter TIME_STEP 					= 32'h27101D7D,							// 2fs time step
	// The home cell this unit is working on
	parameter CELL_X						= 4'd2,
	parameter CELL_Y						= 4'd2,
	parameter CELL_Z						= 4'd2,
	// High level parameters
	parameter NUM_EVAL_UNIT					= 1,									// # of evaluation units in the design
	// Dataset defined parameters
	parameter MAX_CELL_COUNT_PER_DIM 		= 5,									// Maximum cell count among the 3 dimensions
	parameter NUM_NEIGHBOR_CELLS			= 13,									// # of neighbor cells per home cell, for Half-shell method, is 13
	parameter CELL_ID_WIDTH					= 3,									// log(NUM_NEIGHBOR_CELLS)
	parameter MAX_CELL_PARTICLE_NUM			= 290,									// The maximum # of particles can be in a cell
	parameter CELL_ADDR_WIDTH				= 9,									// log(MAX_CELL_PARTICLE_NUM)
	parameter PARTICLE_ID_WIDTH				= CELL_ID_WIDTH*3+CELL_ADDR_WIDTH,		// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	// Filter parameters
	parameter NUM_FILTER					= 8,	//4
	parameter ARBITER_MSB 					= 128,	//8								// 2^(NUM_FILTER-1)
	parameter FILTER_BUFFER_DEPTH 			= 32,
	parameter FILTER_BUFFER_ADDR_WIDTH		= 5,
	parameter CUTOFF_2 						= 32'h43100000,							// (12^2=144 in IEEE floating point)
	// Force Evaluation parameters
	parameter SEGMENT_NUM					= 14,
	parameter SEGMENT_WIDTH					= 4,
	parameter BIN_NUM						= 256,
	parameter BIN_WIDTH						= 8,
	parameter LOOKUP_NUM					= SEGMENT_NUM * BIN_NUM,				// SEGMENT_NUM * BIN_NUM
	parameter LOOKUP_ADDR_WIDTH				= SEGMENT_WIDTH + BIN_WIDTH,			// log LOOKUP_NUM / log 2
	// Force (accmulation) cache parameters
	parameter FORCE_CACHE_BUFFER_DEPTH		= 16,									// Force cache input buffer depth, for partial force accumulation
	parameter FORCE_CACHE_BUFFER_ADDR_WIDTH	= 4										// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
)
(
	input clk,
	input rst,
	input start,
	// These are all temp output ports	output [NUM_EVAL_UNIT*PARTICLE_ID_WIDTH-1:0] ref_particle_id,
	output [NUM_EVAL_UNIT*DATA_WIDTH-1:0] ref_LJ_Force_X,
	output [NUM_EVAL_UNIT*DATA_WIDTH-1:0] ref_LJ_Force_Y,
	output [NUM_EVAL_UNIT*DATA_WIDTH-1:0] ref_LJ_Force_Z,
	output [NUM_EVAL_UNIT-1:0] ref_forceoutput_valid,
	output [NUM_EVAL_UNIT*PARTICLE_ID_WIDTH-1:0] neighbor_particle_id,
	output [NUM_EVAL_UNIT*DATA_WIDTH-1:0] neighbor_LJ_Force_X,
	output [NUM_EVAL_UNIT*DATA_WIDTH-1:0] neighbor_LJ_Force_Y,
	output [NUM_EVAL_UNIT*DATA_WIDTH-1:0] neighbor_LJ_Force_Z,
	output [NUM_EVAL_UNIT-1:0] neighbor_forceoutput_valid,
	// Done signals
	// When entire home cell is done processing, this will keep high until the next time 'start' signal turn high
	output out_home_cell_evaluation_done,
	// When motion update is done processing, remain high until the next motion update starts
	output out_motion_update_done,
	// Dummy signal selecting which cell is the home cell
	// Need a logic to replace this, generate by out_Motion_Update_cur_cell
	input [7:0] in_sel,
	// Dummy output for motion update
	output [3*CELL_ID_WIDTH-1:0] out_Motion_Update_cur_cell
);

	///////////////////////////////////////////////////////////////////////////////////////////////
	// Signals between Cell Module and FSM
	///////////////////////////////////////////////////////////////////////////////////////////////
	//// Signals connect from cell module to FSM
	// Position Data
	// Order: MSB->LSB {333,332,331,323,322,321,313,312,311,233,232,231,223,222} Homecell is on LSB side
	wire [252*3*DATA_WIDTH-1:0] Position_Cache_readout_position;
	//// Signals connect from FSM to cell modules
	wire FSM_to_Cell_rden;
	// Read Address to cells
	wire [CELL_ADDR_WIDTH-1:0] FSM_to_Cell_read_addr;


	///////////////////////////////////////////////////////////////////////////////////////////////
	// Signals between Force Evaluation Unit and Particle Pairs Generation
	///////////////////////////////////////////////////////////////////////////////////////////////
	//// Signals connect from FSM to Force Evaluation module
	wire [NUM_FILTER*3*DATA_WIDTH-1:0] FSM_to_ForceEval_ref_particle_position;
	wire [NUM_FILTER*3*DATA_WIDTH-1:0] FSM_to_ForceEval_neighbor_particle_position;
	wire [NUM_FILTER*PARTICLE_ID_WIDTH-1:0] FSM_to_ForceEval_ref_particle_id;			// {cell_x, cell_y, cell_z, ref_particle_rd_addr}
	wire [NUM_FILTER*PARTICLE_ID_WIDTH-1:0] FSM_to_ForceEval_neighbor_particle_id;		// {cell_x, cell_y, cell_z, neighbor_particle_rd_addr}
	wire [NUM_FILTER-1:0] FSM_to_ForceEval_input_pair_valid;			// Signify the valid of input particle data, this signal should have 1 cycle delay of the rden signal, thus wait for the data read out from BRAM
	//// Signals connect from Force Evaluation module to FSM
	wire [NUM_FILTER-1:0] ForceEval_to_FSM_backpressure;
	wire ForceEval_to_FSM_all_buffer_empty;
	//// Signals handles the reference output valid
	// Special signal to handle the output valid for the last reference particle
	wire FSM_almost_done_generation;
	// Signal connect to the output of Force evaluation valid
	wire ForceEval_ref_output_valid;
	// Generate the 'ref_forceoutput_valid' signal
	assign ref_forceoutput_valid = ForceEval_ref_output_valid || FSM_almost_done_generation;
	

	///////////////////////////////////////////////////////////////////////////////////////////////
	// Motion Update Signals
	///////////////////////////////////////////////////////////////////////////////////////////////
	// Use this signal to locate the rising edge of out_home_cell_evaluation_done signal
	// only start motion update when rising edge is detected
	reg prev_out_home_cell_evaluation_done;
	always@(posedge clk)
		begin
		prev_out_home_cell_evaluation_done <= out_home_cell_evaluation_done;
	end
	wire Motion_Update_start;
	assign Motion_Update_start = (out_home_cell_evaluation_done && prev_out_home_cell_evaluation_done == 0);
	// The enable singal from Motion Update module, this signal will remain high during the entire motion update process
	wire Motion_Update_enable;
	wire [3*CELL_ID_WIDTH-1:0] Motion_Update_cur_cell;
	// Motion Update read in data from caches
	wire [CELL_ADDR_WIDTH-1:0] Motion_Update_position_read_addr;
	wire Motion_Update_position_read_en;
	reg [3*DATA_WIDTH-1:0] Motion_Update_position_data;
	wire [CELL_ADDR_WIDTH-1:0] Motion_Update_force_read_addr;
	wire Motion_Update_force_read_en;
	reg [3*DATA_WIDTH-1:0] Motion_Update_force_data;
	wire [CELL_ADDR_WIDTH-1:0] Motion_Update_velocity_read_addr;
	wire Motion_Update_velocity_read_en;
	reg [3*DATA_WIDTH-1:0] Motion_Update_velocity_data;
	// Motion Update write back data
	wire [3*CELL_ID_WIDTH-1:0] Motion_Update_dst_cell;
	wire [3*DATA_WIDTH-1:0] Motion_Update_out_velocity_data;
	wire Motion_Update_out_velocity_data_valid;
	wire [3*DATA_WIDTH-1:0] Motion_Update_out_position_data;
	wire Motion_Update_out_position_data_valid;
	// Motion Update select input from force caches
	reg [251:0] wire_motion_update_to_cache_read_force_request;
	wire [251:0] wire_cache_to_motion_update_partial_force_valid;
	wire [252*3*DATA_WIDTH-1:0] wire_cache_to_motion_update_partial_force;
	wire [252*PARTICLE_ID_WIDTH-1:0] wire_cache_to_motion_update_particle_id;
	wire [252*3*DATA_WIDTH-1:0] wire_cache_to_motion_update_velocity_data;
	always@(*)
		begin
		wire_motion_update_to_cache_read_force_request <= Motion_Update_enable << in_sel;
		case(in_sel)
			0:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH];
				end
			1:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH];
				end
			2:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH];
				end
			3:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH];
				end
			4:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH];
				end
			5:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH];
				end
			6:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH];
				end
			7:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH];
				end
			8:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[9*3*DATA_WIDTH-1:8*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[9*3*DATA_WIDTH-1:8*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[9*3*DATA_WIDTH-1:8*3*DATA_WIDTH];
				end
			9:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[10*3*DATA_WIDTH-1:9*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[10*3*DATA_WIDTH-1:9*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[10*3*DATA_WIDTH-1:9*3*DATA_WIDTH];
				end
			10:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[11*3*DATA_WIDTH-1:10*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[11*3*DATA_WIDTH-1:10*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[11*3*DATA_WIDTH-1:10*3*DATA_WIDTH];
				end
			11:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[12*3*DATA_WIDTH-1:11*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[12*3*DATA_WIDTH-1:11*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[12*3*DATA_WIDTH-1:11*3*DATA_WIDTH];
				end
			12:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[13*3*DATA_WIDTH-1:12*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[13*3*DATA_WIDTH-1:12*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[13*3*DATA_WIDTH-1:12*3*DATA_WIDTH];
				end
			13:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[14*3*DATA_WIDTH-1:13*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[14*3*DATA_WIDTH-1:13*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[14*3*DATA_WIDTH-1:13*3*DATA_WIDTH];
				end
			14:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[15*3*DATA_WIDTH-1:14*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[15*3*DATA_WIDTH-1:14*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[15*3*DATA_WIDTH-1:14*3*DATA_WIDTH];
				end
			15:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[16*3*DATA_WIDTH-1:15*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[16*3*DATA_WIDTH-1:15*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[16*3*DATA_WIDTH-1:15*3*DATA_WIDTH];
				end
			16:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH];
				end
			17:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH];
				end
			18:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH];
				end
			19:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH];
				end
			20:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH];
				end
			21:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH];
				end
			22:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH];
				end
			23:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH];
				end
			24:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[25*3*DATA_WIDTH-1:24*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[25*3*DATA_WIDTH-1:24*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[25*3*DATA_WIDTH-1:24*3*DATA_WIDTH];
				end
			25:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[26*3*DATA_WIDTH-1:25*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[26*3*DATA_WIDTH-1:25*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[26*3*DATA_WIDTH-1:25*3*DATA_WIDTH];
				end
			26:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[27*3*DATA_WIDTH-1:26*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[27*3*DATA_WIDTH-1:26*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[27*3*DATA_WIDTH-1:26*3*DATA_WIDTH];
				end
			27:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[28*3*DATA_WIDTH-1:27*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[28*3*DATA_WIDTH-1:27*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[28*3*DATA_WIDTH-1:27*3*DATA_WIDTH];
				end
			28:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH];
				end
			29:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH];
				end
			30:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH];
				end
			31:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH];
				end
			32:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[33*3*DATA_WIDTH-1:32*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[33*3*DATA_WIDTH-1:32*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[33*3*DATA_WIDTH-1:32*3*DATA_WIDTH];
				end
			33:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[34*3*DATA_WIDTH-1:33*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[34*3*DATA_WIDTH-1:33*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[34*3*DATA_WIDTH-1:33*3*DATA_WIDTH];
				end
			34:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[35*3*DATA_WIDTH-1:34*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[35*3*DATA_WIDTH-1:34*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[35*3*DATA_WIDTH-1:34*3*DATA_WIDTH];
				end
			35:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[36*3*DATA_WIDTH-1:35*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[36*3*DATA_WIDTH-1:35*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[36*3*DATA_WIDTH-1:35*3*DATA_WIDTH];
				end
			36:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[37*3*DATA_WIDTH-1:36*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[37*3*DATA_WIDTH-1:36*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[37*3*DATA_WIDTH-1:36*3*DATA_WIDTH];
				end
			37:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[38*3*DATA_WIDTH-1:37*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[38*3*DATA_WIDTH-1:37*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[38*3*DATA_WIDTH-1:37*3*DATA_WIDTH];
				end
			38:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[39*3*DATA_WIDTH-1:38*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[39*3*DATA_WIDTH-1:38*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[39*3*DATA_WIDTH-1:38*3*DATA_WIDTH];
				end
			39:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[40*3*DATA_WIDTH-1:39*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[40*3*DATA_WIDTH-1:39*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[40*3*DATA_WIDTH-1:39*3*DATA_WIDTH];
				end
			40:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[41*3*DATA_WIDTH-1:40*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[41*3*DATA_WIDTH-1:40*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[41*3*DATA_WIDTH-1:40*3*DATA_WIDTH];
				end
			41:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[42*3*DATA_WIDTH-1:41*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[42*3*DATA_WIDTH-1:41*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[42*3*DATA_WIDTH-1:41*3*DATA_WIDTH];
				end
			42:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[43*3*DATA_WIDTH-1:42*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[43*3*DATA_WIDTH-1:42*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[43*3*DATA_WIDTH-1:42*3*DATA_WIDTH];
				end
			43:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[44*3*DATA_WIDTH-1:43*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[44*3*DATA_WIDTH-1:43*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[44*3*DATA_WIDTH-1:43*3*DATA_WIDTH];
				end
			44:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[45*3*DATA_WIDTH-1:44*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[45*3*DATA_WIDTH-1:44*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[45*3*DATA_WIDTH-1:44*3*DATA_WIDTH];
				end
			45:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[46*3*DATA_WIDTH-1:45*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[46*3*DATA_WIDTH-1:45*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[46*3*DATA_WIDTH-1:45*3*DATA_WIDTH];
				end
			46:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[47*3*DATA_WIDTH-1:46*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[47*3*DATA_WIDTH-1:46*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[47*3*DATA_WIDTH-1:46*3*DATA_WIDTH];
				end
			47:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[48*3*DATA_WIDTH-1:47*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[48*3*DATA_WIDTH-1:47*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[48*3*DATA_WIDTH-1:47*3*DATA_WIDTH];
				end
			48:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[49*3*DATA_WIDTH-1:48*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[49*3*DATA_WIDTH-1:48*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[49*3*DATA_WIDTH-1:48*3*DATA_WIDTH];
				end
			49:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[50*3*DATA_WIDTH-1:49*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[50*3*DATA_WIDTH-1:49*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[50*3*DATA_WIDTH-1:49*3*DATA_WIDTH];
				end
			50:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[51*3*DATA_WIDTH-1:50*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[51*3*DATA_WIDTH-1:50*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[51*3*DATA_WIDTH-1:50*3*DATA_WIDTH];
				end
			51:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[52*3*DATA_WIDTH-1:51*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[52*3*DATA_WIDTH-1:51*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[52*3*DATA_WIDTH-1:51*3*DATA_WIDTH];
				end
			52:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[53*3*DATA_WIDTH-1:52*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[53*3*DATA_WIDTH-1:52*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[53*3*DATA_WIDTH-1:52*3*DATA_WIDTH];
				end
			53:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[54*3*DATA_WIDTH-1:53*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[54*3*DATA_WIDTH-1:53*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[54*3*DATA_WIDTH-1:53*3*DATA_WIDTH];
				end
			54:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[55*3*DATA_WIDTH-1:54*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[55*3*DATA_WIDTH-1:54*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[55*3*DATA_WIDTH-1:54*3*DATA_WIDTH];
				end
			55:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[56*3*DATA_WIDTH-1:55*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[56*3*DATA_WIDTH-1:55*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[56*3*DATA_WIDTH-1:55*3*DATA_WIDTH];
				end
			56:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[57*3*DATA_WIDTH-1:56*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[57*3*DATA_WIDTH-1:56*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[57*3*DATA_WIDTH-1:56*3*DATA_WIDTH];
				end
			57:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[58*3*DATA_WIDTH-1:57*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[58*3*DATA_WIDTH-1:57*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[58*3*DATA_WIDTH-1:57*3*DATA_WIDTH];
				end
			58:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[59*3*DATA_WIDTH-1:58*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[59*3*DATA_WIDTH-1:58*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[59*3*DATA_WIDTH-1:58*3*DATA_WIDTH];
				end
			59:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[60*3*DATA_WIDTH-1:59*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[60*3*DATA_WIDTH-1:59*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[60*3*DATA_WIDTH-1:59*3*DATA_WIDTH];
				end
			60:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[61*3*DATA_WIDTH-1:60*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[61*3*DATA_WIDTH-1:60*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[61*3*DATA_WIDTH-1:60*3*DATA_WIDTH];
				end
			61:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[62*3*DATA_WIDTH-1:61*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[62*3*DATA_WIDTH-1:61*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[62*3*DATA_WIDTH-1:61*3*DATA_WIDTH];
				end
			62:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[63*3*DATA_WIDTH-1:62*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[63*3*DATA_WIDTH-1:62*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[63*3*DATA_WIDTH-1:62*3*DATA_WIDTH];
				end
			63:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[64*3*DATA_WIDTH-1:63*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[64*3*DATA_WIDTH-1:63*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[64*3*DATA_WIDTH-1:63*3*DATA_WIDTH];
				end
			64:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[65*3*DATA_WIDTH-1:64*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[65*3*DATA_WIDTH-1:64*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[65*3*DATA_WIDTH-1:64*3*DATA_WIDTH];
				end
			65:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[66*3*DATA_WIDTH-1:65*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[66*3*DATA_WIDTH-1:65*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[66*3*DATA_WIDTH-1:65*3*DATA_WIDTH];
				end
			66:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[67*3*DATA_WIDTH-1:66*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[67*3*DATA_WIDTH-1:66*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[67*3*DATA_WIDTH-1:66*3*DATA_WIDTH];
				end
			67:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[68*3*DATA_WIDTH-1:67*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[68*3*DATA_WIDTH-1:67*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[68*3*DATA_WIDTH-1:67*3*DATA_WIDTH];
				end
			68:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[69*3*DATA_WIDTH-1:68*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[69*3*DATA_WIDTH-1:68*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[69*3*DATA_WIDTH-1:68*3*DATA_WIDTH];
				end
			69:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[70*3*DATA_WIDTH-1:69*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[70*3*DATA_WIDTH-1:69*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[70*3*DATA_WIDTH-1:69*3*DATA_WIDTH];
				end
			70:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[71*3*DATA_WIDTH-1:70*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[71*3*DATA_WIDTH-1:70*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[71*3*DATA_WIDTH-1:70*3*DATA_WIDTH];
				end
			71:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[72*3*DATA_WIDTH-1:71*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[72*3*DATA_WIDTH-1:71*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[72*3*DATA_WIDTH-1:71*3*DATA_WIDTH];
				end
			72:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[73*3*DATA_WIDTH-1:72*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[73*3*DATA_WIDTH-1:72*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[73*3*DATA_WIDTH-1:72*3*DATA_WIDTH];
				end
			73:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[74*3*DATA_WIDTH-1:73*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[74*3*DATA_WIDTH-1:73*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[74*3*DATA_WIDTH-1:73*3*DATA_WIDTH];
				end
			74:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[75*3*DATA_WIDTH-1:74*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[75*3*DATA_WIDTH-1:74*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[75*3*DATA_WIDTH-1:74*3*DATA_WIDTH];
				end
			75:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[76*3*DATA_WIDTH-1:75*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[76*3*DATA_WIDTH-1:75*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[76*3*DATA_WIDTH-1:75*3*DATA_WIDTH];
				end
			76:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[77*3*DATA_WIDTH-1:76*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[77*3*DATA_WIDTH-1:76*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[77*3*DATA_WIDTH-1:76*3*DATA_WIDTH];
				end
			77:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[78*3*DATA_WIDTH-1:77*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[78*3*DATA_WIDTH-1:77*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[78*3*DATA_WIDTH-1:77*3*DATA_WIDTH];
				end
			78:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[79*3*DATA_WIDTH-1:78*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[79*3*DATA_WIDTH-1:78*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[79*3*DATA_WIDTH-1:78*3*DATA_WIDTH];
				end
			79:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[80*3*DATA_WIDTH-1:79*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[80*3*DATA_WIDTH-1:79*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[80*3*DATA_WIDTH-1:79*3*DATA_WIDTH];
				end
			80:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[81*3*DATA_WIDTH-1:80*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[81*3*DATA_WIDTH-1:80*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[81*3*DATA_WIDTH-1:80*3*DATA_WIDTH];
				end
			81:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[82*3*DATA_WIDTH-1:81*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[82*3*DATA_WIDTH-1:81*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[82*3*DATA_WIDTH-1:81*3*DATA_WIDTH];
				end
			82:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[83*3*DATA_WIDTH-1:82*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[83*3*DATA_WIDTH-1:82*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[83*3*DATA_WIDTH-1:82*3*DATA_WIDTH];
				end
			83:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[84*3*DATA_WIDTH-1:83*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[84*3*DATA_WIDTH-1:83*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[84*3*DATA_WIDTH-1:83*3*DATA_WIDTH];
				end
			84:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[85*3*DATA_WIDTH-1:84*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[85*3*DATA_WIDTH-1:84*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[85*3*DATA_WIDTH-1:84*3*DATA_WIDTH];
				end
			85:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[86*3*DATA_WIDTH-1:85*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[86*3*DATA_WIDTH-1:85*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[86*3*DATA_WIDTH-1:85*3*DATA_WIDTH];
				end
			86:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[87*3*DATA_WIDTH-1:86*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[87*3*DATA_WIDTH-1:86*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[87*3*DATA_WIDTH-1:86*3*DATA_WIDTH];
				end
			87:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[88*3*DATA_WIDTH-1:87*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[88*3*DATA_WIDTH-1:87*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[88*3*DATA_WIDTH-1:87*3*DATA_WIDTH];
				end
			88:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[89*3*DATA_WIDTH-1:88*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[89*3*DATA_WIDTH-1:88*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[89*3*DATA_WIDTH-1:88*3*DATA_WIDTH];
				end
			89:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[90*3*DATA_WIDTH-1:89*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[90*3*DATA_WIDTH-1:89*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[90*3*DATA_WIDTH-1:89*3*DATA_WIDTH];
				end
			90:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[91*3*DATA_WIDTH-1:90*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[91*3*DATA_WIDTH-1:90*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[91*3*DATA_WIDTH-1:90*3*DATA_WIDTH];
				end
			91:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[92*3*DATA_WIDTH-1:91*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[92*3*DATA_WIDTH-1:91*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[92*3*DATA_WIDTH-1:91*3*DATA_WIDTH];
				end
			92:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[93*3*DATA_WIDTH-1:92*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[93*3*DATA_WIDTH-1:92*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[93*3*DATA_WIDTH-1:92*3*DATA_WIDTH];
				end
			93:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[94*3*DATA_WIDTH-1:93*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[94*3*DATA_WIDTH-1:93*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[94*3*DATA_WIDTH-1:93*3*DATA_WIDTH];
				end
			94:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[95*3*DATA_WIDTH-1:94*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[95*3*DATA_WIDTH-1:94*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[95*3*DATA_WIDTH-1:94*3*DATA_WIDTH];
				end
			95:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[96*3*DATA_WIDTH-1:95*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[96*3*DATA_WIDTH-1:95*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[96*3*DATA_WIDTH-1:95*3*DATA_WIDTH];
				end
			96:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[97*3*DATA_WIDTH-1:96*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[97*3*DATA_WIDTH-1:96*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[97*3*DATA_WIDTH-1:96*3*DATA_WIDTH];
				end
			97:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[98*3*DATA_WIDTH-1:97*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[98*3*DATA_WIDTH-1:97*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[98*3*DATA_WIDTH-1:97*3*DATA_WIDTH];
				end
			98:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[99*3*DATA_WIDTH-1:98*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[99*3*DATA_WIDTH-1:98*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[99*3*DATA_WIDTH-1:98*3*DATA_WIDTH];
				end
			99:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[100*3*DATA_WIDTH-1:99*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[100*3*DATA_WIDTH-1:99*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[100*3*DATA_WIDTH-1:99*3*DATA_WIDTH];
				end
			100:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[101*3*DATA_WIDTH-1:100*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[101*3*DATA_WIDTH-1:100*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[101*3*DATA_WIDTH-1:100*3*DATA_WIDTH];
				end
			101:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[102*3*DATA_WIDTH-1:101*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[102*3*DATA_WIDTH-1:101*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[102*3*DATA_WIDTH-1:101*3*DATA_WIDTH];
				end
			102:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[103*3*DATA_WIDTH-1:102*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[103*3*DATA_WIDTH-1:102*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[103*3*DATA_WIDTH-1:102*3*DATA_WIDTH];
				end
			103:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[104*3*DATA_WIDTH-1:103*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[104*3*DATA_WIDTH-1:103*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[104*3*DATA_WIDTH-1:103*3*DATA_WIDTH];
				end
			104:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[105*3*DATA_WIDTH-1:104*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[105*3*DATA_WIDTH-1:104*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[105*3*DATA_WIDTH-1:104*3*DATA_WIDTH];
				end
			105:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[106*3*DATA_WIDTH-1:105*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[106*3*DATA_WIDTH-1:105*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[106*3*DATA_WIDTH-1:105*3*DATA_WIDTH];
				end
			106:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[107*3*DATA_WIDTH-1:106*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[107*3*DATA_WIDTH-1:106*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[107*3*DATA_WIDTH-1:106*3*DATA_WIDTH];
				end
			107:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[108*3*DATA_WIDTH-1:107*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[108*3*DATA_WIDTH-1:107*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[108*3*DATA_WIDTH-1:107*3*DATA_WIDTH];
				end
			108:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[109*3*DATA_WIDTH-1:108*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[109*3*DATA_WIDTH-1:108*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[109*3*DATA_WIDTH-1:108*3*DATA_WIDTH];
				end
			109:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[110*3*DATA_WIDTH-1:109*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[110*3*DATA_WIDTH-1:109*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[110*3*DATA_WIDTH-1:109*3*DATA_WIDTH];
				end
			110:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[111*3*DATA_WIDTH-1:110*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[111*3*DATA_WIDTH-1:110*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[111*3*DATA_WIDTH-1:110*3*DATA_WIDTH];
				end
			111:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[112*3*DATA_WIDTH-1:111*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[112*3*DATA_WIDTH-1:111*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[112*3*DATA_WIDTH-1:111*3*DATA_WIDTH];
				end
			112:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[113*3*DATA_WIDTH-1:112*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[113*3*DATA_WIDTH-1:112*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[113*3*DATA_WIDTH-1:112*3*DATA_WIDTH];
				end
			113:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[114*3*DATA_WIDTH-1:113*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[114*3*DATA_WIDTH-1:113*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[114*3*DATA_WIDTH-1:113*3*DATA_WIDTH];
				end
			114:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[115*3*DATA_WIDTH-1:114*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[115*3*DATA_WIDTH-1:114*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[115*3*DATA_WIDTH-1:114*3*DATA_WIDTH];
				end
			115:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[116*3*DATA_WIDTH-1:115*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[116*3*DATA_WIDTH-1:115*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[116*3*DATA_WIDTH-1:115*3*DATA_WIDTH];
				end
			116:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[117*3*DATA_WIDTH-1:116*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[117*3*DATA_WIDTH-1:116*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[117*3*DATA_WIDTH-1:116*3*DATA_WIDTH];
				end
			117:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[118*3*DATA_WIDTH-1:117*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[118*3*DATA_WIDTH-1:117*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[118*3*DATA_WIDTH-1:117*3*DATA_WIDTH];
				end
			118:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[119*3*DATA_WIDTH-1:118*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[119*3*DATA_WIDTH-1:118*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[119*3*DATA_WIDTH-1:118*3*DATA_WIDTH];
				end
			119:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[120*3*DATA_WIDTH-1:119*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[120*3*DATA_WIDTH-1:119*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[120*3*DATA_WIDTH-1:119*3*DATA_WIDTH];
				end
			120:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[121*3*DATA_WIDTH-1:120*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[121*3*DATA_WIDTH-1:120*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[121*3*DATA_WIDTH-1:120*3*DATA_WIDTH];
				end
			121:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[122*3*DATA_WIDTH-1:121*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[122*3*DATA_WIDTH-1:121*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[122*3*DATA_WIDTH-1:121*3*DATA_WIDTH];
				end
			122:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[123*3*DATA_WIDTH-1:122*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[123*3*DATA_WIDTH-1:122*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[123*3*DATA_WIDTH-1:122*3*DATA_WIDTH];
				end
			123:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[124*3*DATA_WIDTH-1:123*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[124*3*DATA_WIDTH-1:123*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[124*3*DATA_WIDTH-1:123*3*DATA_WIDTH];
				end
			124:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[125*3*DATA_WIDTH-1:124*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[125*3*DATA_WIDTH-1:124*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[125*3*DATA_WIDTH-1:124*3*DATA_WIDTH];
				end
			125:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[126*3*DATA_WIDTH-1:125*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[126*3*DATA_WIDTH-1:125*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[126*3*DATA_WIDTH-1:125*3*DATA_WIDTH];
				end
			126:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[127*3*DATA_WIDTH-1:126*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[127*3*DATA_WIDTH-1:126*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[127*3*DATA_WIDTH-1:126*3*DATA_WIDTH];
				end
			127:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[128*3*DATA_WIDTH-1:127*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[128*3*DATA_WIDTH-1:127*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[128*3*DATA_WIDTH-1:127*3*DATA_WIDTH];
				end
			128:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[129*3*DATA_WIDTH-1:128*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[129*3*DATA_WIDTH-1:128*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[129*3*DATA_WIDTH-1:128*3*DATA_WIDTH];
				end
			129:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[130*3*DATA_WIDTH-1:129*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[130*3*DATA_WIDTH-1:129*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[130*3*DATA_WIDTH-1:129*3*DATA_WIDTH];
				end
			130:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[131*3*DATA_WIDTH-1:130*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[131*3*DATA_WIDTH-1:130*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[131*3*DATA_WIDTH-1:130*3*DATA_WIDTH];
				end
			131:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[132*3*DATA_WIDTH-1:131*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[132*3*DATA_WIDTH-1:131*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[132*3*DATA_WIDTH-1:131*3*DATA_WIDTH];
				end
			132:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[133*3*DATA_WIDTH-1:132*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[133*3*DATA_WIDTH-1:132*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[133*3*DATA_WIDTH-1:132*3*DATA_WIDTH];
				end
			133:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[134*3*DATA_WIDTH-1:133*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[134*3*DATA_WIDTH-1:133*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[134*3*DATA_WIDTH-1:133*3*DATA_WIDTH];
				end
			134:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[135*3*DATA_WIDTH-1:134*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[135*3*DATA_WIDTH-1:134*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[135*3*DATA_WIDTH-1:134*3*DATA_WIDTH];
				end
			135:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[136*3*DATA_WIDTH-1:135*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[136*3*DATA_WIDTH-1:135*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[136*3*DATA_WIDTH-1:135*3*DATA_WIDTH];
				end
			136:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[137*3*DATA_WIDTH-1:136*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[137*3*DATA_WIDTH-1:136*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[137*3*DATA_WIDTH-1:136*3*DATA_WIDTH];
				end
			137:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[138*3*DATA_WIDTH-1:137*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[138*3*DATA_WIDTH-1:137*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[138*3*DATA_WIDTH-1:137*3*DATA_WIDTH];
				end
			138:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[139*3*DATA_WIDTH-1:138*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[139*3*DATA_WIDTH-1:138*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[139*3*DATA_WIDTH-1:138*3*DATA_WIDTH];
				end
			139:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[140*3*DATA_WIDTH-1:139*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[140*3*DATA_WIDTH-1:139*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[140*3*DATA_WIDTH-1:139*3*DATA_WIDTH];
				end
			140:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[141*3*DATA_WIDTH-1:140*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[141*3*DATA_WIDTH-1:140*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[141*3*DATA_WIDTH-1:140*3*DATA_WIDTH];
				end
			141:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[142*3*DATA_WIDTH-1:141*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[142*3*DATA_WIDTH-1:141*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[142*3*DATA_WIDTH-1:141*3*DATA_WIDTH];
				end
			142:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[143*3*DATA_WIDTH-1:142*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[143*3*DATA_WIDTH-1:142*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[143*3*DATA_WIDTH-1:142*3*DATA_WIDTH];
				end
			143:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[144*3*DATA_WIDTH-1:143*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[144*3*DATA_WIDTH-1:143*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[144*3*DATA_WIDTH-1:143*3*DATA_WIDTH];
				end
			144:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[145*3*DATA_WIDTH-1:144*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[145*3*DATA_WIDTH-1:144*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[145*3*DATA_WIDTH-1:144*3*DATA_WIDTH];
				end
			145:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[146*3*DATA_WIDTH-1:145*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[146*3*DATA_WIDTH-1:145*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[146*3*DATA_WIDTH-1:145*3*DATA_WIDTH];
				end
			146:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[147*3*DATA_WIDTH-1:146*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[147*3*DATA_WIDTH-1:146*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[147*3*DATA_WIDTH-1:146*3*DATA_WIDTH];
				end
			147:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[148*3*DATA_WIDTH-1:147*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[148*3*DATA_WIDTH-1:147*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[148*3*DATA_WIDTH-1:147*3*DATA_WIDTH];
				end
			148:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[149*3*DATA_WIDTH-1:148*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[149*3*DATA_WIDTH-1:148*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[149*3*DATA_WIDTH-1:148*3*DATA_WIDTH];
				end
			149:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[150*3*DATA_WIDTH-1:149*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[150*3*DATA_WIDTH-1:149*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[150*3*DATA_WIDTH-1:149*3*DATA_WIDTH];
				end
			150:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[151*3*DATA_WIDTH-1:150*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[151*3*DATA_WIDTH-1:150*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[151*3*DATA_WIDTH-1:150*3*DATA_WIDTH];
				end
			151:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[152*3*DATA_WIDTH-1:151*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[152*3*DATA_WIDTH-1:151*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[152*3*DATA_WIDTH-1:151*3*DATA_WIDTH];
				end
			152:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[153*3*DATA_WIDTH-1:152*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[153*3*DATA_WIDTH-1:152*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[153*3*DATA_WIDTH-1:152*3*DATA_WIDTH];
				end
			153:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[154*3*DATA_WIDTH-1:153*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[154*3*DATA_WIDTH-1:153*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[154*3*DATA_WIDTH-1:153*3*DATA_WIDTH];
				end
			154:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[155*3*DATA_WIDTH-1:154*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[155*3*DATA_WIDTH-1:154*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[155*3*DATA_WIDTH-1:154*3*DATA_WIDTH];
				end
			155:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[156*3*DATA_WIDTH-1:155*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[156*3*DATA_WIDTH-1:155*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[156*3*DATA_WIDTH-1:155*3*DATA_WIDTH];
				end
			156:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[157*3*DATA_WIDTH-1:156*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[157*3*DATA_WIDTH-1:156*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[157*3*DATA_WIDTH-1:156*3*DATA_WIDTH];
				end
			157:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[158*3*DATA_WIDTH-1:157*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[158*3*DATA_WIDTH-1:157*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[158*3*DATA_WIDTH-1:157*3*DATA_WIDTH];
				end
			158:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[159*3*DATA_WIDTH-1:158*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[159*3*DATA_WIDTH-1:158*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[159*3*DATA_WIDTH-1:158*3*DATA_WIDTH];
				end
			159:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[160*3*DATA_WIDTH-1:159*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[160*3*DATA_WIDTH-1:159*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[160*3*DATA_WIDTH-1:159*3*DATA_WIDTH];
				end
			160:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[161*3*DATA_WIDTH-1:160*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[161*3*DATA_WIDTH-1:160*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[161*3*DATA_WIDTH-1:160*3*DATA_WIDTH];
				end
			161:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[162*3*DATA_WIDTH-1:161*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[162*3*DATA_WIDTH-1:161*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[162*3*DATA_WIDTH-1:161*3*DATA_WIDTH];
				end
			162:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[163*3*DATA_WIDTH-1:162*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[163*3*DATA_WIDTH-1:162*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[163*3*DATA_WIDTH-1:162*3*DATA_WIDTH];
				end
			163:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[164*3*DATA_WIDTH-1:163*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[164*3*DATA_WIDTH-1:163*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[164*3*DATA_WIDTH-1:163*3*DATA_WIDTH];
				end
			164:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[165*3*DATA_WIDTH-1:164*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[165*3*DATA_WIDTH-1:164*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[165*3*DATA_WIDTH-1:164*3*DATA_WIDTH];
				end
			165:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[166*3*DATA_WIDTH-1:165*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[166*3*DATA_WIDTH-1:165*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[166*3*DATA_WIDTH-1:165*3*DATA_WIDTH];
				end
			166:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[167*3*DATA_WIDTH-1:166*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[167*3*DATA_WIDTH-1:166*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[167*3*DATA_WIDTH-1:166*3*DATA_WIDTH];
				end
			167:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[168*3*DATA_WIDTH-1:167*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[168*3*DATA_WIDTH-1:167*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[168*3*DATA_WIDTH-1:167*3*DATA_WIDTH];
				end
			168:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[169*3*DATA_WIDTH-1:168*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[169*3*DATA_WIDTH-1:168*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[169*3*DATA_WIDTH-1:168*3*DATA_WIDTH];
				end
			169:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[170*3*DATA_WIDTH-1:169*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[170*3*DATA_WIDTH-1:169*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[170*3*DATA_WIDTH-1:169*3*DATA_WIDTH];
				end
			170:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[171*3*DATA_WIDTH-1:170*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[171*3*DATA_WIDTH-1:170*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[171*3*DATA_WIDTH-1:170*3*DATA_WIDTH];
				end
			171:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[172*3*DATA_WIDTH-1:171*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[172*3*DATA_WIDTH-1:171*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[172*3*DATA_WIDTH-1:171*3*DATA_WIDTH];
				end
			172:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[173*3*DATA_WIDTH-1:172*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[173*3*DATA_WIDTH-1:172*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[173*3*DATA_WIDTH-1:172*3*DATA_WIDTH];
				end
			173:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[174*3*DATA_WIDTH-1:173*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[174*3*DATA_WIDTH-1:173*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[174*3*DATA_WIDTH-1:173*3*DATA_WIDTH];
				end
			174:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[175*3*DATA_WIDTH-1:174*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[175*3*DATA_WIDTH-1:174*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[175*3*DATA_WIDTH-1:174*3*DATA_WIDTH];
				end
			175:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[176*3*DATA_WIDTH-1:175*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[176*3*DATA_WIDTH-1:175*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[176*3*DATA_WIDTH-1:175*3*DATA_WIDTH];
				end
			176:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[177*3*DATA_WIDTH-1:176*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[177*3*DATA_WIDTH-1:176*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[177*3*DATA_WIDTH-1:176*3*DATA_WIDTH];
				end
			177:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[178*3*DATA_WIDTH-1:177*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[178*3*DATA_WIDTH-1:177*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[178*3*DATA_WIDTH-1:177*3*DATA_WIDTH];
				end
			178:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[179*3*DATA_WIDTH-1:178*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[179*3*DATA_WIDTH-1:178*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[179*3*DATA_WIDTH-1:178*3*DATA_WIDTH];
				end
			179:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[180*3*DATA_WIDTH-1:179*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[180*3*DATA_WIDTH-1:179*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[180*3*DATA_WIDTH-1:179*3*DATA_WIDTH];
				end
			180:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[181*3*DATA_WIDTH-1:180*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[181*3*DATA_WIDTH-1:180*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[181*3*DATA_WIDTH-1:180*3*DATA_WIDTH];
				end
			181:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[182*3*DATA_WIDTH-1:181*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[182*3*DATA_WIDTH-1:181*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[182*3*DATA_WIDTH-1:181*3*DATA_WIDTH];
				end
			182:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[183*3*DATA_WIDTH-1:182*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[183*3*DATA_WIDTH-1:182*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[183*3*DATA_WIDTH-1:182*3*DATA_WIDTH];
				end
			183:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[184*3*DATA_WIDTH-1:183*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[184*3*DATA_WIDTH-1:183*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[184*3*DATA_WIDTH-1:183*3*DATA_WIDTH];
				end
			184:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[185*3*DATA_WIDTH-1:184*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[185*3*DATA_WIDTH-1:184*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[185*3*DATA_WIDTH-1:184*3*DATA_WIDTH];
				end
			185:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[186*3*DATA_WIDTH-1:185*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[186*3*DATA_WIDTH-1:185*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[186*3*DATA_WIDTH-1:185*3*DATA_WIDTH];
				end
			186:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[187*3*DATA_WIDTH-1:186*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[187*3*DATA_WIDTH-1:186*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[187*3*DATA_WIDTH-1:186*3*DATA_WIDTH];
				end
			187:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[188*3*DATA_WIDTH-1:187*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[188*3*DATA_WIDTH-1:187*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[188*3*DATA_WIDTH-1:187*3*DATA_WIDTH];
				end
			188:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[189*3*DATA_WIDTH-1:188*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[189*3*DATA_WIDTH-1:188*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[189*3*DATA_WIDTH-1:188*3*DATA_WIDTH];
				end
			189:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[190*3*DATA_WIDTH-1:189*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[190*3*DATA_WIDTH-1:189*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[190*3*DATA_WIDTH-1:189*3*DATA_WIDTH];
				end
			190:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[191*3*DATA_WIDTH-1:190*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[191*3*DATA_WIDTH-1:190*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[191*3*DATA_WIDTH-1:190*3*DATA_WIDTH];
				end
			191:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[192*3*DATA_WIDTH-1:191*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[192*3*DATA_WIDTH-1:191*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[192*3*DATA_WIDTH-1:191*3*DATA_WIDTH];
				end
			192:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[193*3*DATA_WIDTH-1:192*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[193*3*DATA_WIDTH-1:192*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[193*3*DATA_WIDTH-1:192*3*DATA_WIDTH];
				end
			193:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[194*3*DATA_WIDTH-1:193*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[194*3*DATA_WIDTH-1:193*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[194*3*DATA_WIDTH-1:193*3*DATA_WIDTH];
				end
			194:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[195*3*DATA_WIDTH-1:194*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[195*3*DATA_WIDTH-1:194*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[195*3*DATA_WIDTH-1:194*3*DATA_WIDTH];
				end
			195:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[196*3*DATA_WIDTH-1:195*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[196*3*DATA_WIDTH-1:195*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[196*3*DATA_WIDTH-1:195*3*DATA_WIDTH];
				end
			196:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[197*3*DATA_WIDTH-1:196*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[197*3*DATA_WIDTH-1:196*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[197*3*DATA_WIDTH-1:196*3*DATA_WIDTH];
				end
			197:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[198*3*DATA_WIDTH-1:197*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[198*3*DATA_WIDTH-1:197*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[198*3*DATA_WIDTH-1:197*3*DATA_WIDTH];
				end
			198:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[199*3*DATA_WIDTH-1:198*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[199*3*DATA_WIDTH-1:198*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[199*3*DATA_WIDTH-1:198*3*DATA_WIDTH];
				end
			199:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[200*3*DATA_WIDTH-1:199*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[200*3*DATA_WIDTH-1:199*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[200*3*DATA_WIDTH-1:199*3*DATA_WIDTH];
				end
			200:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[201*3*DATA_WIDTH-1:200*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[201*3*DATA_WIDTH-1:200*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[201*3*DATA_WIDTH-1:200*3*DATA_WIDTH];
				end
			201:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[202*3*DATA_WIDTH-1:201*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[202*3*DATA_WIDTH-1:201*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[202*3*DATA_WIDTH-1:201*3*DATA_WIDTH];
				end
			202:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[203*3*DATA_WIDTH-1:202*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[203*3*DATA_WIDTH-1:202*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[203*3*DATA_WIDTH-1:202*3*DATA_WIDTH];
				end
			203:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[204*3*DATA_WIDTH-1:203*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[204*3*DATA_WIDTH-1:203*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[204*3*DATA_WIDTH-1:203*3*DATA_WIDTH];
				end
			204:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[205*3*DATA_WIDTH-1:204*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[205*3*DATA_WIDTH-1:204*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[205*3*DATA_WIDTH-1:204*3*DATA_WIDTH];
				end
			205:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[206*3*DATA_WIDTH-1:205*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[206*3*DATA_WIDTH-1:205*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[206*3*DATA_WIDTH-1:205*3*DATA_WIDTH];
				end
			206:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[207*3*DATA_WIDTH-1:206*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[207*3*DATA_WIDTH-1:206*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[207*3*DATA_WIDTH-1:206*3*DATA_WIDTH];
				end
			207:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[208*3*DATA_WIDTH-1:207*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[208*3*DATA_WIDTH-1:207*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[208*3*DATA_WIDTH-1:207*3*DATA_WIDTH];
				end
			208:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[209*3*DATA_WIDTH-1:208*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[209*3*DATA_WIDTH-1:208*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[209*3*DATA_WIDTH-1:208*3*DATA_WIDTH];
				end
			209:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[210*3*DATA_WIDTH-1:209*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[210*3*DATA_WIDTH-1:209*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[210*3*DATA_WIDTH-1:209*3*DATA_WIDTH];
				end
			210:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[211*3*DATA_WIDTH-1:210*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[211*3*DATA_WIDTH-1:210*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[211*3*DATA_WIDTH-1:210*3*DATA_WIDTH];
				end
			211:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[212*3*DATA_WIDTH-1:211*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[212*3*DATA_WIDTH-1:211*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[212*3*DATA_WIDTH-1:211*3*DATA_WIDTH];
				end
			212:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[213*3*DATA_WIDTH-1:212*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[213*3*DATA_WIDTH-1:212*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[213*3*DATA_WIDTH-1:212*3*DATA_WIDTH];
				end
			213:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[214*3*DATA_WIDTH-1:213*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[214*3*DATA_WIDTH-1:213*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[214*3*DATA_WIDTH-1:213*3*DATA_WIDTH];
				end
			214:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[215*3*DATA_WIDTH-1:214*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[215*3*DATA_WIDTH-1:214*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[215*3*DATA_WIDTH-1:214*3*DATA_WIDTH];
				end
			215:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[216*3*DATA_WIDTH-1:215*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[216*3*DATA_WIDTH-1:215*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[216*3*DATA_WIDTH-1:215*3*DATA_WIDTH];
				end
			216:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[217*3*DATA_WIDTH-1:216*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[217*3*DATA_WIDTH-1:216*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[217*3*DATA_WIDTH-1:216*3*DATA_WIDTH];
				end
			217:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[218*3*DATA_WIDTH-1:217*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[218*3*DATA_WIDTH-1:217*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[218*3*DATA_WIDTH-1:217*3*DATA_WIDTH];
				end
			218:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[219*3*DATA_WIDTH-1:218*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[219*3*DATA_WIDTH-1:218*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[219*3*DATA_WIDTH-1:218*3*DATA_WIDTH];
				end
			219:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[220*3*DATA_WIDTH-1:219*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[220*3*DATA_WIDTH-1:219*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[220*3*DATA_WIDTH-1:219*3*DATA_WIDTH];
				end
			220:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[221*3*DATA_WIDTH-1:220*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[221*3*DATA_WIDTH-1:220*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[221*3*DATA_WIDTH-1:220*3*DATA_WIDTH];
				end
			221:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[222*3*DATA_WIDTH-1:221*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[222*3*DATA_WIDTH-1:221*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[222*3*DATA_WIDTH-1:221*3*DATA_WIDTH];
				end
			222:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[223*3*DATA_WIDTH-1:222*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[223*3*DATA_WIDTH-1:222*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[223*3*DATA_WIDTH-1:222*3*DATA_WIDTH];
				end
			223:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[224*3*DATA_WIDTH-1:223*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[224*3*DATA_WIDTH-1:223*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[224*3*DATA_WIDTH-1:223*3*DATA_WIDTH];
				end
			224:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[225*3*DATA_WIDTH-1:224*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[225*3*DATA_WIDTH-1:224*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[225*3*DATA_WIDTH-1:224*3*DATA_WIDTH];
				end
			225:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[226*3*DATA_WIDTH-1:225*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[226*3*DATA_WIDTH-1:225*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[226*3*DATA_WIDTH-1:225*3*DATA_WIDTH];
				end
			226:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[227*3*DATA_WIDTH-1:226*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[227*3*DATA_WIDTH-1:226*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[227*3*DATA_WIDTH-1:226*3*DATA_WIDTH];
				end
			227:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[228*3*DATA_WIDTH-1:227*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[228*3*DATA_WIDTH-1:227*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[228*3*DATA_WIDTH-1:227*3*DATA_WIDTH];
				end
			228:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[229*3*DATA_WIDTH-1:228*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[229*3*DATA_WIDTH-1:228*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[229*3*DATA_WIDTH-1:228*3*DATA_WIDTH];
				end
			229:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[230*3*DATA_WIDTH-1:229*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[230*3*DATA_WIDTH-1:229*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[230*3*DATA_WIDTH-1:229*3*DATA_WIDTH];
				end
			230:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[231*3*DATA_WIDTH-1:230*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[231*3*DATA_WIDTH-1:230*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[231*3*DATA_WIDTH-1:230*3*DATA_WIDTH];
				end
			231:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[232*3*DATA_WIDTH-1:231*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[232*3*DATA_WIDTH-1:231*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[232*3*DATA_WIDTH-1:231*3*DATA_WIDTH];
				end
			232:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[233*3*DATA_WIDTH-1:232*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[233*3*DATA_WIDTH-1:232*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[233*3*DATA_WIDTH-1:232*3*DATA_WIDTH];
				end
			233:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[234*3*DATA_WIDTH-1:233*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[234*3*DATA_WIDTH-1:233*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[234*3*DATA_WIDTH-1:233*3*DATA_WIDTH];
				end
			234:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[235*3*DATA_WIDTH-1:234*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[235*3*DATA_WIDTH-1:234*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[235*3*DATA_WIDTH-1:234*3*DATA_WIDTH];
				end
			235:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[236*3*DATA_WIDTH-1:235*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[236*3*DATA_WIDTH-1:235*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[236*3*DATA_WIDTH-1:235*3*DATA_WIDTH];
				end
			236:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[237*3*DATA_WIDTH-1:236*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[237*3*DATA_WIDTH-1:236*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[237*3*DATA_WIDTH-1:236*3*DATA_WIDTH];
				end
			237:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[238*3*DATA_WIDTH-1:237*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[238*3*DATA_WIDTH-1:237*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[238*3*DATA_WIDTH-1:237*3*DATA_WIDTH];
				end
			238:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[239*3*DATA_WIDTH-1:238*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[239*3*DATA_WIDTH-1:238*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[239*3*DATA_WIDTH-1:238*3*DATA_WIDTH];
				end
			239:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[240*3*DATA_WIDTH-1:239*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[240*3*DATA_WIDTH-1:239*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[240*3*DATA_WIDTH-1:239*3*DATA_WIDTH];
				end
			240:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[241*3*DATA_WIDTH-1:240*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[241*3*DATA_WIDTH-1:240*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[241*3*DATA_WIDTH-1:240*3*DATA_WIDTH];
				end
			241:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[242*3*DATA_WIDTH-1:241*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[242*3*DATA_WIDTH-1:241*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[242*3*DATA_WIDTH-1:241*3*DATA_WIDTH];
				end
			242:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[243*3*DATA_WIDTH-1:242*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[243*3*DATA_WIDTH-1:242*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[243*3*DATA_WIDTH-1:242*3*DATA_WIDTH];
				end
			243:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[244*3*DATA_WIDTH-1:243*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[244*3*DATA_WIDTH-1:243*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[244*3*DATA_WIDTH-1:243*3*DATA_WIDTH];
				end
			244:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[245*3*DATA_WIDTH-1:244*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[245*3*DATA_WIDTH-1:244*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[245*3*DATA_WIDTH-1:244*3*DATA_WIDTH];
				end
			245:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[246*3*DATA_WIDTH-1:245*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[246*3*DATA_WIDTH-1:245*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[246*3*DATA_WIDTH-1:245*3*DATA_WIDTH];
				end
			246:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[247*3*DATA_WIDTH-1:246*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[247*3*DATA_WIDTH-1:246*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[247*3*DATA_WIDTH-1:246*3*DATA_WIDTH];
				end
			247:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[248*3*DATA_WIDTH-1:247*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[248*3*DATA_WIDTH-1:247*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[248*3*DATA_WIDTH-1:247*3*DATA_WIDTH];
				end
			248:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[249*3*DATA_WIDTH-1:248*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[249*3*DATA_WIDTH-1:248*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[249*3*DATA_WIDTH-1:248*3*DATA_WIDTH];
				end
			249:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[250*3*DATA_WIDTH-1:249*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[250*3*DATA_WIDTH-1:249*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[250*3*DATA_WIDTH-1:249*3*DATA_WIDTH];
				end
			250:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[251*3*DATA_WIDTH-1:250*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[251*3*DATA_WIDTH-1:250*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[251*3*DATA_WIDTH-1:250*3*DATA_WIDTH];
				end
			251:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[252*3*DATA_WIDTH-1:251*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[252*3*DATA_WIDTH-1:251*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[252*3*DATA_WIDTH-1:251*3*DATA_WIDTH];
				end
			default:
				begin
				Motion_Update_position_data <= Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH];
				Motion_Update_force_data <= wire_cache_to_motion_update_partial_force[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH];
				Motion_Update_velocity_data <= wire_cache_to_motion_update_velocity_data[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH];
				end
		endcase
		end


	///////////////////////////////////////////////////////////////////////////////////////////////
	// FSM for generating particle pairs
	///////////////////////////////////////////////////////////////////////////////////////////////
	Particle_Pair_Gen_Dummy
	#(
		.DATA_WIDTH(DATA_WIDTH),
		// The # of cells in each dimension
		.CELL_X_NUM(7),
		.CELL_Y_NUM(7),
		.CELL_Z_NUM(7),
		.TOTAL_CELL_NUM(252),
		// High level parameters
		.NUM_EVAL_UNIT(NUM_EVAL_UNIT),							// # of evaluation units in the design
		// Dataset defined parameters
		.NUM_NEIGHBOR_CELLS(NUM_NEIGHBOR_CELLS),				// # of neighbor cells per home cell, for Half-shell method, is 13
		.CELL_ID_WIDTH(CELL_ID_WIDTH),							// log(NUM_NEIGHBOR_CELLS)
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),						// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH),					// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		// Filter parameters
		.NUM_FILTER(NUM_FILTER),
		.ARBITER_MSB(ARBITER_MSB),									// 2^(NUM_FILTER-1)
		.FILTER_BUFFER_DEPTH(FILTER_BUFFER_DEPTH),
		.FILTER_BUFFER_ADDR_WIDTH(FILTER_BUFFER_ADDR_WIDTH)
	)
	Particle_Pair_Gen
	(
		.clk(clk),
		.rst(rst),
		.start(start),
		// Ports connect to Cell Memory Module
		// Order: MSB->LSB {333,332,331,323,322,321,313,312,311,233,232,231,223,222} Homecell is on LSB side
		.Cell_to_FSM_readout_particle_position(Position_Cache_readout_position),					// input  [(NUM_NEIGHBOR_CELLS+1)*3*DATA_WIDTH-1:0] 
		.FSM_to_Cell_read_addr(FSM_to_Cell_read_addr),																// output [(NUM_NEIGHBOR_CELLS+1)*CELL_ADDR_WIDTH-1:0] 
		.FSM_to_Cell_rden(FSM_to_Cell_rden),
		// Ports connect to Force Evaluation Unit
		.ForceEval_to_FSM_backpressure(ForceEval_to_FSM_backpressure),											// input  [NUM_FILTER-1:0]  								// Backpressure signal from Force Evaluation Unit
		.ForceEval_to_FSM_all_buffer_empty(ForceEval_to_FSM_all_buffer_empty),								// input															// Only when all the filter buffers are empty, then the FSM will move on to the next reference particle
		.FSM_to_ForceEval_ref_particle_position(FSM_to_ForceEval_ref_particle_position),  				// output [NUM_FILTER*3*DATA_WIDTH-1:0] 
		.FSM_to_ForceEval_neighbor_particle_position(FSM_to_ForceEval_neighbor_particle_position),	// output [NUM_FILTER*3*DATA_WIDTH-1:0] 
		.FSM_to_ForceEval_ref_particle_id(FSM_to_ForceEval_ref_particle_id),									// output [NUM_FILTER*PARTICLE_ID_WIDTH-1:0] 		// {cell_z, cell_y, cell_x, ref_particle_rd_addr}
		.FSM_to_ForceEval_neighbor_particle_id(FSM_to_ForceEval_neighbor_particle_id),					// output [NUM_FILTER*PARTICLE_ID_WIDTH-1:0] 		// {cell_z, cell_y, cell_x, neighbor_particle_rd_addr}
		.FSM_to_ForceEval_input_pair_valid(FSM_to_ForceEval_input_pair_valid),								// output reg [NUM_FILTER-1:0]   						// Signify the valid of input particle data, this signal should have 1 cycle delay of the rden signal, thus wait for the data read out from BRAM
		// Special signal to handle the output valid for the last reference particle
		.FSM_almost_done_generation(FSM_almost_done_generation),
		// Ports to top level modules
		.done(out_home_cell_evaluation_done)
	);


	///////////////////////////////////////////////////////////////////////////////////////////////
	// Force evaluation and accumulation unit
	///////////////////////////////////////////////////////////////////////////////////////////////
	RL_LJ_Evaluation_Unit
	#(
		.DATA_WIDTH(DATA_WIDTH),
		// The home cell this unit is working on (Not been used so far)
		.CELL_X(CELL_X),
		.CELL_Y(CELL_Y),
		.CELL_Z(CELL_Z),
		// Dataset defined parameters
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH),
		// Filter parameters
		.NUM_FILTER(NUM_FILTER),
		.ARBITER_MSB(ARBITER_MSB),
		.FILTER_BUFFER_DEPTH(FILTER_BUFFER_DEPTH),
		.FILTER_BUFFER_ADDR_WIDTH(FILTER_BUFFER_ADDR_WIDTH),
		.CUTOFF_2(CUTOFF_2),
		// Force Evaluation parameters
		.SEGMENT_NUM(SEGMENT_NUM),
		.SEGMENT_WIDTH(SEGMENT_WIDTH),
		.BIN_NUM(BIN_NUM),
		.BIN_WIDTH(BIN_WIDTH),
		.LOOKUP_NUM(LOOKUP_NUM),
		.LOOKUP_ADDR_WIDTH(LOOKUP_ADDR_WIDTH)
	)
	RL_LJ_Evaluation_Unit
	(
		.clk(clk),
		.rst(rst),
		.in_input_pair_valid(FSM_to_ForceEval_input_pair_valid),						//input  [NUM_FILTER-1:0]
		.in_ref_particle_id(FSM_to_ForceEval_ref_particle_id),							//input  [NUM_FILTER*PARTICLE_ID_WIDTH-1:0]
		.in_neighbor_particle_id(FSM_to_ForceEval_neighbor_particle_id),				//input  [NUM_FILTER*PARTICLE_ID_WIDTH-1:0]
		.in_ref_particle_position(FSM_to_ForceEval_ref_particle_position),				//input  [NUM_FILTER*3*DATA_WIDTH-1:0]			// {refz, refy, refx}
		.in_neighbor_particle_position(FSM_to_ForceEval_neighbor_particle_position),	//input  [NUM_FILTER*3*DATA_WIDTH-1:0]			// {neighborz, neighbory, neighborx}
		.out_back_pressure_to_input(ForceEval_to_FSM_backpressure),					//output [NUM_FILTER-1:0] 						// backpressure signal to stop new data arrival from particle memory
		.out_all_buffer_empty_to_input(ForceEval_to_FSM_all_buffer_empty),				//output										// Only when all the filter buffers are empty, then the FSM will move on to the next reference particle
		// Output accumulated force for reference particles
		// The output value is the accumulated value
		// Connected to home cell
		.out_ref_particle_id(ref_particle_id),						//output [PARTICLE_ID_WIDTH-1:0]
		.out_ref_LJ_Force_X(ref_LJ_Force_X),						//output [DATA_WIDTH-1:0]
		.out_ref_LJ_Force_Y(ref_LJ_Force_Y),						//output [DATA_WIDTH-1:0]
		.out_ref_LJ_Force_Z(ref_LJ_Force_Z),						//output [DATA_WIDTH-1:0]
		.out_ref_force_valid(ForceEval_ref_output_valid),			//output
		// Output partial force for neighbor particles
		// The output value should be the minus value of the calculated force data
		// Connected to neighbor cells, if the neighbor paritle comes from the home cell, then discard, since the value will be recalculated when evaluating this particle as reference one
		.out_neighbor_particle_id(neighbor_particle_id),			//output [PARTICLE_ID_WIDTH-1:0]
		.out_neighbor_LJ_Force_X(neighbor_LJ_Force_X),				//output [DATA_WIDTH-1:0]
		.out_neighbor_LJ_Force_Y(neighbor_LJ_Force_Y),				//output [DATA_WIDTH-1:0]
		.out_neighbor_LJ_Force_Z(neighbor_LJ_Force_Z),				//output [DATA_WIDTH-1:0]
		.out_neighbor_force_valid(neighbor_forceoutput_valid)		//output
	);

	///////////////////////////////////////////////////////////////////////////////////////////////
	// Motion Update Unit
	// This Unit can work on multiple cells, or a single cell
	///////////////////////////////////////////////////////////////////////////////////////////////
	// Assign output signal
	assign out_Motion_Update_cur_cell = Motion_Update_cur_cell;
	Motion_Update
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.TIME_STEP(TIME_STEP),										// 2fs time step
		// Cell id this unit related to
		.CELL_X(CELL_X),
		.CELL_Y(CELL_Y),
		.CELL_Z(CELL_Z),
		// Dataset defined parameters
		.MAX_CELL_COUNT_PER_DIM(MAX_CELL_COUNT_PER_DIM),			// Maximum cell count among the 3 dimensions
		.CELL_ID_WIDTH(CELL_ID_WIDTH),								// log(NUM_NEIGHBOR_CELLS)
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),				// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),							// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)						// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	)
	Motion_Update
	(
		.clk(clk),
		.rst(rst),
		.motion_update_start(Motion_Update_start),					// Start Motion update after the home cell is done evaluating
		.motion_update_done(out_motion_update_done),					// Remain high until the next motion update starts
		// Output the targeting home cell
		// When this module is responsible for multiple cells, then the control signal is broadcast to multiple cells, while a mux need to implement on the input side to select from those cells
		.out_cur_working_cell_x(Motion_Update_cur_cell[3*CELL_ID_WIDTH-1:2*CELL_ID_WIDTH]),
		.out_cur_working_cell_y(Motion_Update_cur_cell[2*CELL_ID_WIDTH-1:1*CELL_ID_WIDTH]),
		.out_cur_working_cell_z(Motion_Update_cur_cell[1*CELL_ID_WIDTH-1:0*CELL_ID_WIDTH]),
		// Read from Position Cache
		.in_position_data(Motion_Update_position_data),
		.out_position_cache_rd_en(Motion_Update_position_read_en),
		.out_position_cache_rd_addr(Motion_Update_position_read_addr),
		// Read from Force Cache
		.in_force_data(Motion_Update_force_data),
		.out_force_cache_rd_en(Motion_Update_force_read_en),
		.out_force_cache_rd_addr(Motion_Update_force_read_addr),
		// Read from Velocity Cache
		.in_velocity_data(Motion_Update_velocity_data),
		.out_velocity_cache_rd_en(Motion_Update_velocity_read_en),
		.out_velocity_cache_rd_addr(Motion_Update_velocity_read_addr),
		// Motion update enable signal
		.out_motion_update_enable(Motion_Update_enable),		// Remine high during the entire motion update process
		// Write back to Velocity Cache
		.out_velocity_data(Motion_Update_out_velocity_data),	// The updated velocity value
		.out_velocity_data_valid(Motion_Update_out_velocity_data_valid),
		.out_velocity_destination_cell(Motion_Update_dst_cell),
		// Write back to Position Cache
		.out_position_data(Motion_Update_out_position_data),
		.out_position_data_valid(Motion_Update_out_position_data_valid),
		.out_position_destination_cell()						// Leave this one idle, the value is the same as out_velocity_destination_cell
	);

	///////////////////////////////////////////////////////////////////////////////////////////////
	// Cell particle memory
	// In this impelementation, take cell(2,2,2) as home cell for example (cell cooridinate starts from (1,1,1))
	// The neighbor cells including:
	// Side: (3,1,1),(3,1,2),(3,1,3),(3,2,1),(3,2,2),(3,2,3),(3,3,1),(3,3,2),(3,3,3)
	// Column: (2,3,1),(2,3,2),(2,3,3)
	// Top: (2,2,3)
	// Data orgainization in cell memory: (pos_z, pos_y, pos_x)
	///////////////////////////////////////////////////////////////////////////////////////////////
	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(1)
	)
	Pos_Cache_1_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(2)
	)
	Pos_Cache_1_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(3)
	)
	Pos_Cache_1_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(4)
	)
	Pos_Cache_1_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(5)
	)
	Pos_Cache_1_1_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(6)
	)
	Pos_Cache_1_1_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(1)
	)
	Pos_Cache_1_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(2)
	)
	Pos_Cache_1_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(3)
	)
	Pos_Cache_1_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[9*3*DATA_WIDTH-1:8*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(4)
	)
	Pos_Cache_1_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[10*3*DATA_WIDTH-1:9*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(5)
	)
	Pos_Cache_1_2_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[11*3*DATA_WIDTH-1:10*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(6)
	)
	Pos_Cache_1_2_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[12*3*DATA_WIDTH-1:11*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(1)
	)
	Pos_Cache_1_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[13*3*DATA_WIDTH-1:12*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(2)
	)
	Pos_Cache_1_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[14*3*DATA_WIDTH-1:13*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(3)
	)
	Pos_Cache_1_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[15*3*DATA_WIDTH-1:14*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(4)
	)
	Pos_Cache_1_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[16*3*DATA_WIDTH-1:15*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(5)
	)
	Pos_Cache_1_3_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(6)
	)
	Pos_Cache_1_3_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(1)
	)
	Pos_Cache_1_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(2)
	)
	Pos_Cache_1_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(3)
	)
	Pos_Cache_1_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(4)
	)
	Pos_Cache_1_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(5)
	)
	Pos_Cache_1_4_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(6)
	)
	Pos_Cache_1_4_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(5),
		.CELL_Z(1)
	)
	Pos_Cache_1_5_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[25*3*DATA_WIDTH-1:24*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(5),
		.CELL_Z(2)
	)
	Pos_Cache_1_5_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[26*3*DATA_WIDTH-1:25*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(5),
		.CELL_Z(3)
	)
	Pos_Cache_1_5_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[27*3*DATA_WIDTH-1:26*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(5),
		.CELL_Z(4)
	)
	Pos_Cache_1_5_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[28*3*DATA_WIDTH-1:27*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(5),
		.CELL_Z(5)
	)
	Pos_Cache_1_5_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(5),
		.CELL_Z(6)
	)
	Pos_Cache_1_5_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(6),
		.CELL_Z(1)
	)
	Pos_Cache_1_6_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(6),
		.CELL_Z(2)
	)
	Pos_Cache_1_6_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(6),
		.CELL_Z(3)
	)
	Pos_Cache_1_6_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[33*3*DATA_WIDTH-1:32*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(6),
		.CELL_Z(4)
	)
	Pos_Cache_1_6_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[34*3*DATA_WIDTH-1:33*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(6),
		.CELL_Z(5)
	)
	Pos_Cache_1_6_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[35*3*DATA_WIDTH-1:34*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(6),
		.CELL_Z(6)
	)
	Pos_Cache_1_6_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[36*3*DATA_WIDTH-1:35*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(1)
	)
	Pos_Cache_2_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[37*3*DATA_WIDTH-1:36*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(2)
	)
	Pos_Cache_2_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[38*3*DATA_WIDTH-1:37*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(3)
	)
	Pos_Cache_2_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[39*3*DATA_WIDTH-1:38*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(4)
	)
	Pos_Cache_2_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[40*3*DATA_WIDTH-1:39*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(5)
	)
	Pos_Cache_2_1_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[41*3*DATA_WIDTH-1:40*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(6)
	)
	Pos_Cache_2_1_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[42*3*DATA_WIDTH-1:41*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(1)
	)
	Pos_Cache_2_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[43*3*DATA_WIDTH-1:42*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(2)
	)
	Pos_Cache_2_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[44*3*DATA_WIDTH-1:43*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(3)
	)
	Pos_Cache_2_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[45*3*DATA_WIDTH-1:44*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(4)
	)
	Pos_Cache_2_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[46*3*DATA_WIDTH-1:45*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(5)
	)
	Pos_Cache_2_2_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[47*3*DATA_WIDTH-1:46*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(6)
	)
	Pos_Cache_2_2_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[48*3*DATA_WIDTH-1:47*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(1)
	)
	Pos_Cache_2_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[49*3*DATA_WIDTH-1:48*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(2)
	)
	Pos_Cache_2_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[50*3*DATA_WIDTH-1:49*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(3)
	)
	Pos_Cache_2_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[51*3*DATA_WIDTH-1:50*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(4)
	)
	Pos_Cache_2_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[52*3*DATA_WIDTH-1:51*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(5)
	)
	Pos_Cache_2_3_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[53*3*DATA_WIDTH-1:52*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(6)
	)
	Pos_Cache_2_3_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[54*3*DATA_WIDTH-1:53*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(1)
	)
	Pos_Cache_2_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[55*3*DATA_WIDTH-1:54*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(2)
	)
	Pos_Cache_2_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[56*3*DATA_WIDTH-1:55*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(3)
	)
	Pos_Cache_2_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[57*3*DATA_WIDTH-1:56*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(4)
	)
	Pos_Cache_2_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[58*3*DATA_WIDTH-1:57*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(5)
	)
	Pos_Cache_2_4_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[59*3*DATA_WIDTH-1:58*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(6)
	)
	Pos_Cache_2_4_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[60*3*DATA_WIDTH-1:59*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(5),
		.CELL_Z(1)
	)
	Pos_Cache_2_5_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[61*3*DATA_WIDTH-1:60*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(5),
		.CELL_Z(2)
	)
	Pos_Cache_2_5_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[62*3*DATA_WIDTH-1:61*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(5),
		.CELL_Z(3)
	)
	Pos_Cache_2_5_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[63*3*DATA_WIDTH-1:62*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(5),
		.CELL_Z(4)
	)
	Pos_Cache_2_5_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[64*3*DATA_WIDTH-1:63*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(5),
		.CELL_Z(5)
	)
	Pos_Cache_2_5_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[65*3*DATA_WIDTH-1:64*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(5),
		.CELL_Z(6)
	)
	Pos_Cache_2_5_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[66*3*DATA_WIDTH-1:65*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(6),
		.CELL_Z(1)
	)
	Pos_Cache_2_6_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[67*3*DATA_WIDTH-1:66*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(6),
		.CELL_Z(2)
	)
	Pos_Cache_2_6_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[68*3*DATA_WIDTH-1:67*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(6),
		.CELL_Z(3)
	)
	Pos_Cache_2_6_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[69*3*DATA_WIDTH-1:68*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(6),
		.CELL_Z(4)
	)
	Pos_Cache_2_6_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[70*3*DATA_WIDTH-1:69*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(6),
		.CELL_Z(5)
	)
	Pos_Cache_2_6_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[71*3*DATA_WIDTH-1:70*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(6),
		.CELL_Z(6)
	)
	Pos_Cache_2_6_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[72*3*DATA_WIDTH-1:71*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(1)
	)
	Pos_Cache_3_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[73*3*DATA_WIDTH-1:72*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(2)
	)
	Pos_Cache_3_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[74*3*DATA_WIDTH-1:73*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(3)
	)
	Pos_Cache_3_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[75*3*DATA_WIDTH-1:74*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(4)
	)
	Pos_Cache_3_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[76*3*DATA_WIDTH-1:75*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(5)
	)
	Pos_Cache_3_1_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[77*3*DATA_WIDTH-1:76*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(6)
	)
	Pos_Cache_3_1_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[78*3*DATA_WIDTH-1:77*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(1)
	)
	Pos_Cache_3_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[79*3*DATA_WIDTH-1:78*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(2)
	)
	Pos_Cache_3_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[80*3*DATA_WIDTH-1:79*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(3)
	)
	Pos_Cache_3_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[81*3*DATA_WIDTH-1:80*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(4)
	)
	Pos_Cache_3_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[82*3*DATA_WIDTH-1:81*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(5)
	)
	Pos_Cache_3_2_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[83*3*DATA_WIDTH-1:82*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(6)
	)
	Pos_Cache_3_2_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[84*3*DATA_WIDTH-1:83*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(1)
	)
	Pos_Cache_3_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[85*3*DATA_WIDTH-1:84*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(2)
	)
	Pos_Cache_3_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[86*3*DATA_WIDTH-1:85*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(3)
	)
	Pos_Cache_3_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[87*3*DATA_WIDTH-1:86*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(4)
	)
	Pos_Cache_3_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[88*3*DATA_WIDTH-1:87*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(5)
	)
	Pos_Cache_3_3_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[89*3*DATA_WIDTH-1:88*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(6)
	)
	Pos_Cache_3_3_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[90*3*DATA_WIDTH-1:89*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(1)
	)
	Pos_Cache_3_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[91*3*DATA_WIDTH-1:90*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(2)
	)
	Pos_Cache_3_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[92*3*DATA_WIDTH-1:91*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(3)
	)
	Pos_Cache_3_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[93*3*DATA_WIDTH-1:92*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(4)
	)
	Pos_Cache_3_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[94*3*DATA_WIDTH-1:93*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(5)
	)
	Pos_Cache_3_4_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[95*3*DATA_WIDTH-1:94*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(6)
	)
	Pos_Cache_3_4_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[96*3*DATA_WIDTH-1:95*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(5),
		.CELL_Z(1)
	)
	Pos_Cache_3_5_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[97*3*DATA_WIDTH-1:96*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(5),
		.CELL_Z(2)
	)
	Pos_Cache_3_5_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[98*3*DATA_WIDTH-1:97*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(5),
		.CELL_Z(3)
	)
	Pos_Cache_3_5_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[99*3*DATA_WIDTH-1:98*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(5),
		.CELL_Z(4)
	)
	Pos_Cache_3_5_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[100*3*DATA_WIDTH-1:99*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(5),
		.CELL_Z(5)
	)
	Pos_Cache_3_5_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[101*3*DATA_WIDTH-1:100*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(5),
		.CELL_Z(6)
	)
	Pos_Cache_3_5_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[102*3*DATA_WIDTH-1:101*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(6),
		.CELL_Z(1)
	)
	Pos_Cache_3_6_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[103*3*DATA_WIDTH-1:102*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(6),
		.CELL_Z(2)
	)
	Pos_Cache_3_6_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[104*3*DATA_WIDTH-1:103*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(6),
		.CELL_Z(3)
	)
	Pos_Cache_3_6_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[105*3*DATA_WIDTH-1:104*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(6),
		.CELL_Z(4)
	)
	Pos_Cache_3_6_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[106*3*DATA_WIDTH-1:105*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(6),
		.CELL_Z(5)
	)
	Pos_Cache_3_6_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[107*3*DATA_WIDTH-1:106*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(6),
		.CELL_Z(6)
	)
	Pos_Cache_3_6_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[108*3*DATA_WIDTH-1:107*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(1)
	)
	Pos_Cache_4_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[109*3*DATA_WIDTH-1:108*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(2)
	)
	Pos_Cache_4_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[110*3*DATA_WIDTH-1:109*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(3)
	)
	Pos_Cache_4_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[111*3*DATA_WIDTH-1:110*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(4)
	)
	Pos_Cache_4_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[112*3*DATA_WIDTH-1:111*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(5)
	)
	Pos_Cache_4_1_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[113*3*DATA_WIDTH-1:112*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(6)
	)
	Pos_Cache_4_1_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[114*3*DATA_WIDTH-1:113*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(1)
	)
	Pos_Cache_4_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[115*3*DATA_WIDTH-1:114*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(2)
	)
	Pos_Cache_4_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[116*3*DATA_WIDTH-1:115*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(3)
	)
	Pos_Cache_4_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[117*3*DATA_WIDTH-1:116*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(4)
	)
	Pos_Cache_4_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[118*3*DATA_WIDTH-1:117*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(5)
	)
	Pos_Cache_4_2_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[119*3*DATA_WIDTH-1:118*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(6)
	)
	Pos_Cache_4_2_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[120*3*DATA_WIDTH-1:119*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(1)
	)
	Pos_Cache_4_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[121*3*DATA_WIDTH-1:120*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(2)
	)
	Pos_Cache_4_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[122*3*DATA_WIDTH-1:121*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(3)
	)
	Pos_Cache_4_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[123*3*DATA_WIDTH-1:122*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(4)
	)
	Pos_Cache_4_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[124*3*DATA_WIDTH-1:123*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(5)
	)
	Pos_Cache_4_3_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[125*3*DATA_WIDTH-1:124*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(6)
	)
	Pos_Cache_4_3_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[126*3*DATA_WIDTH-1:125*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(1)
	)
	Pos_Cache_4_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[127*3*DATA_WIDTH-1:126*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(2)
	)
	Pos_Cache_4_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[128*3*DATA_WIDTH-1:127*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(3)
	)
	Pos_Cache_4_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[129*3*DATA_WIDTH-1:128*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(4)
	)
	Pos_Cache_4_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[130*3*DATA_WIDTH-1:129*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(5)
	)
	Pos_Cache_4_4_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[131*3*DATA_WIDTH-1:130*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(6)
	)
	Pos_Cache_4_4_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[132*3*DATA_WIDTH-1:131*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(5),
		.CELL_Z(1)
	)
	Pos_Cache_4_5_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[133*3*DATA_WIDTH-1:132*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(5),
		.CELL_Z(2)
	)
	Pos_Cache_4_5_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[134*3*DATA_WIDTH-1:133*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(5),
		.CELL_Z(3)
	)
	Pos_Cache_4_5_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[135*3*DATA_WIDTH-1:134*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(5),
		.CELL_Z(4)
	)
	Pos_Cache_4_5_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[136*3*DATA_WIDTH-1:135*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(5),
		.CELL_Z(5)
	)
	Pos_Cache_4_5_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[137*3*DATA_WIDTH-1:136*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(5),
		.CELL_Z(6)
	)
	Pos_Cache_4_5_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[138*3*DATA_WIDTH-1:137*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(6),
		.CELL_Z(1)
	)
	Pos_Cache_4_6_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[139*3*DATA_WIDTH-1:138*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(6),
		.CELL_Z(2)
	)
	Pos_Cache_4_6_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[140*3*DATA_WIDTH-1:139*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(6),
		.CELL_Z(3)
	)
	Pos_Cache_4_6_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[141*3*DATA_WIDTH-1:140*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(6),
		.CELL_Z(4)
	)
	Pos_Cache_4_6_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[142*3*DATA_WIDTH-1:141*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(6),
		.CELL_Z(5)
	)
	Pos_Cache_4_6_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[143*3*DATA_WIDTH-1:142*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(6),
		.CELL_Z(6)
	)
	Pos_Cache_4_6_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[144*3*DATA_WIDTH-1:143*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(1),
		.CELL_Z(1)
	)
	Pos_Cache_5_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[145*3*DATA_WIDTH-1:144*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(1),
		.CELL_Z(2)
	)
	Pos_Cache_5_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[146*3*DATA_WIDTH-1:145*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(1),
		.CELL_Z(3)
	)
	Pos_Cache_5_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[147*3*DATA_WIDTH-1:146*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(1),
		.CELL_Z(4)
	)
	Pos_Cache_5_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[148*3*DATA_WIDTH-1:147*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(1),
		.CELL_Z(5)
	)
	Pos_Cache_5_1_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[149*3*DATA_WIDTH-1:148*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(1),
		.CELL_Z(6)
	)
	Pos_Cache_5_1_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[150*3*DATA_WIDTH-1:149*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(2),
		.CELL_Z(1)
	)
	Pos_Cache_5_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[151*3*DATA_WIDTH-1:150*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(2),
		.CELL_Z(2)
	)
	Pos_Cache_5_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[152*3*DATA_WIDTH-1:151*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(2),
		.CELL_Z(3)
	)
	Pos_Cache_5_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[153*3*DATA_WIDTH-1:152*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(2),
		.CELL_Z(4)
	)
	Pos_Cache_5_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[154*3*DATA_WIDTH-1:153*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(2),
		.CELL_Z(5)
	)
	Pos_Cache_5_2_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[155*3*DATA_WIDTH-1:154*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(2),
		.CELL_Z(6)
	)
	Pos_Cache_5_2_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[156*3*DATA_WIDTH-1:155*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(3),
		.CELL_Z(1)
	)
	Pos_Cache_5_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[157*3*DATA_WIDTH-1:156*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(3),
		.CELL_Z(2)
	)
	Pos_Cache_5_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[158*3*DATA_WIDTH-1:157*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(3),
		.CELL_Z(3)
	)
	Pos_Cache_5_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[159*3*DATA_WIDTH-1:158*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(3),
		.CELL_Z(4)
	)
	Pos_Cache_5_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[160*3*DATA_WIDTH-1:159*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(3),
		.CELL_Z(5)
	)
	Pos_Cache_5_3_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[161*3*DATA_WIDTH-1:160*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(3),
		.CELL_Z(6)
	)
	Pos_Cache_5_3_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[162*3*DATA_WIDTH-1:161*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(4),
		.CELL_Z(1)
	)
	Pos_Cache_5_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[163*3*DATA_WIDTH-1:162*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(4),
		.CELL_Z(2)
	)
	Pos_Cache_5_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[164*3*DATA_WIDTH-1:163*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(4),
		.CELL_Z(3)
	)
	Pos_Cache_5_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[165*3*DATA_WIDTH-1:164*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(4),
		.CELL_Z(4)
	)
	Pos_Cache_5_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[166*3*DATA_WIDTH-1:165*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(4),
		.CELL_Z(5)
	)
	Pos_Cache_5_4_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[167*3*DATA_WIDTH-1:166*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(4),
		.CELL_Z(6)
	)
	Pos_Cache_5_4_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[168*3*DATA_WIDTH-1:167*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(5),
		.CELL_Z(1)
	)
	Pos_Cache_5_5_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[169*3*DATA_WIDTH-1:168*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(5),
		.CELL_Z(2)
	)
	Pos_Cache_5_5_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[170*3*DATA_WIDTH-1:169*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(5),
		.CELL_Z(3)
	)
	Pos_Cache_5_5_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[171*3*DATA_WIDTH-1:170*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(5),
		.CELL_Z(4)
	)
	Pos_Cache_5_5_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[172*3*DATA_WIDTH-1:171*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(5),
		.CELL_Z(5)
	)
	Pos_Cache_5_5_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[173*3*DATA_WIDTH-1:172*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(5),
		.CELL_Z(6)
	)
	Pos_Cache_5_5_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[174*3*DATA_WIDTH-1:173*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(6),
		.CELL_Z(1)
	)
	Pos_Cache_5_6_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[175*3*DATA_WIDTH-1:174*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(6),
		.CELL_Z(2)
	)
	Pos_Cache_5_6_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[176*3*DATA_WIDTH-1:175*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(6),
		.CELL_Z(3)
	)
	Pos_Cache_5_6_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[177*3*DATA_WIDTH-1:176*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(6),
		.CELL_Z(4)
	)
	Pos_Cache_5_6_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[178*3*DATA_WIDTH-1:177*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(6),
		.CELL_Z(5)
	)
	Pos_Cache_5_6_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[179*3*DATA_WIDTH-1:178*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(6),
		.CELL_Z(6)
	)
	Pos_Cache_5_6_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[180*3*DATA_WIDTH-1:179*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(1),
		.CELL_Z(1)
	)
	Pos_Cache_6_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[181*3*DATA_WIDTH-1:180*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(1),
		.CELL_Z(2)
	)
	Pos_Cache_6_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[182*3*DATA_WIDTH-1:181*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(1),
		.CELL_Z(3)
	)
	Pos_Cache_6_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[183*3*DATA_WIDTH-1:182*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(1),
		.CELL_Z(4)
	)
	Pos_Cache_6_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[184*3*DATA_WIDTH-1:183*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(1),
		.CELL_Z(5)
	)
	Pos_Cache_6_1_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[185*3*DATA_WIDTH-1:184*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(1),
		.CELL_Z(6)
	)
	Pos_Cache_6_1_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[186*3*DATA_WIDTH-1:185*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(2),
		.CELL_Z(1)
	)
	Pos_Cache_6_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[187*3*DATA_WIDTH-1:186*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(2),
		.CELL_Z(2)
	)
	Pos_Cache_6_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[188*3*DATA_WIDTH-1:187*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(2),
		.CELL_Z(3)
	)
	Pos_Cache_6_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[189*3*DATA_WIDTH-1:188*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(2),
		.CELL_Z(4)
	)
	Pos_Cache_6_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[190*3*DATA_WIDTH-1:189*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(2),
		.CELL_Z(5)
	)
	Pos_Cache_6_2_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[191*3*DATA_WIDTH-1:190*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(2),
		.CELL_Z(6)
	)
	Pos_Cache_6_2_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[192*3*DATA_WIDTH-1:191*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(3),
		.CELL_Z(1)
	)
	Pos_Cache_6_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[193*3*DATA_WIDTH-1:192*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(3),
		.CELL_Z(2)
	)
	Pos_Cache_6_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[194*3*DATA_WIDTH-1:193*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(3),
		.CELL_Z(3)
	)
	Pos_Cache_6_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[195*3*DATA_WIDTH-1:194*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(3),
		.CELL_Z(4)
	)
	Pos_Cache_6_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[196*3*DATA_WIDTH-1:195*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(3),
		.CELL_Z(5)
	)
	Pos_Cache_6_3_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[197*3*DATA_WIDTH-1:196*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(3),
		.CELL_Z(6)
	)
	Pos_Cache_6_3_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[198*3*DATA_WIDTH-1:197*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(4),
		.CELL_Z(1)
	)
	Pos_Cache_6_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[199*3*DATA_WIDTH-1:198*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(4),
		.CELL_Z(2)
	)
	Pos_Cache_6_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[200*3*DATA_WIDTH-1:199*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(4),
		.CELL_Z(3)
	)
	Pos_Cache_6_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[201*3*DATA_WIDTH-1:200*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(4),
		.CELL_Z(4)
	)
	Pos_Cache_6_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[202*3*DATA_WIDTH-1:201*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(4),
		.CELL_Z(5)
	)
	Pos_Cache_6_4_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[203*3*DATA_WIDTH-1:202*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(4),
		.CELL_Z(6)
	)
	Pos_Cache_6_4_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[204*3*DATA_WIDTH-1:203*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(5),
		.CELL_Z(1)
	)
	Pos_Cache_6_5_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[205*3*DATA_WIDTH-1:204*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(5),
		.CELL_Z(2)
	)
	Pos_Cache_6_5_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[206*3*DATA_WIDTH-1:205*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(5),
		.CELL_Z(3)
	)
	Pos_Cache_6_5_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[207*3*DATA_WIDTH-1:206*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(5),
		.CELL_Z(4)
	)
	Pos_Cache_6_5_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[208*3*DATA_WIDTH-1:207*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(5),
		.CELL_Z(5)
	)
	Pos_Cache_6_5_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[209*3*DATA_WIDTH-1:208*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(5),
		.CELL_Z(6)
	)
	Pos_Cache_6_5_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[210*3*DATA_WIDTH-1:209*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(6),
		.CELL_Z(1)
	)
	Pos_Cache_6_6_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[211*3*DATA_WIDTH-1:210*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(6),
		.CELL_Z(2)
	)
	Pos_Cache_6_6_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[212*3*DATA_WIDTH-1:211*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(6),
		.CELL_Z(3)
	)
	Pos_Cache_6_6_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[213*3*DATA_WIDTH-1:212*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(6),
		.CELL_Z(4)
	)
	Pos_Cache_6_6_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[214*3*DATA_WIDTH-1:213*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(6),
		.CELL_Z(5)
	)
	Pos_Cache_6_6_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[215*3*DATA_WIDTH-1:214*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(6),
		.CELL_Z(6)
	)
	Pos_Cache_6_6_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[216*3*DATA_WIDTH-1:215*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(1),
		.CELL_Z(1)
	)
	Pos_Cache_7_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[217*3*DATA_WIDTH-1:216*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(1),
		.CELL_Z(2)
	)
	Pos_Cache_7_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[218*3*DATA_WIDTH-1:217*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(1),
		.CELL_Z(3)
	)
	Pos_Cache_7_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[219*3*DATA_WIDTH-1:218*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(1),
		.CELL_Z(4)
	)
	Pos_Cache_7_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[220*3*DATA_WIDTH-1:219*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(1),
		.CELL_Z(5)
	)
	Pos_Cache_7_1_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[221*3*DATA_WIDTH-1:220*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(1),
		.CELL_Z(6)
	)
	Pos_Cache_7_1_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[222*3*DATA_WIDTH-1:221*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(2),
		.CELL_Z(1)
	)
	Pos_Cache_7_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[223*3*DATA_WIDTH-1:222*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(2),
		.CELL_Z(2)
	)
	Pos_Cache_7_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[224*3*DATA_WIDTH-1:223*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(2),
		.CELL_Z(3)
	)
	Pos_Cache_7_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[225*3*DATA_WIDTH-1:224*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(2),
		.CELL_Z(4)
	)
	Pos_Cache_7_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[226*3*DATA_WIDTH-1:225*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(2),
		.CELL_Z(5)
	)
	Pos_Cache_7_2_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[227*3*DATA_WIDTH-1:226*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(2),
		.CELL_Z(6)
	)
	Pos_Cache_7_2_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[228*3*DATA_WIDTH-1:227*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(3),
		.CELL_Z(1)
	)
	Pos_Cache_7_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[229*3*DATA_WIDTH-1:228*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(3),
		.CELL_Z(2)
	)
	Pos_Cache_7_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[230*3*DATA_WIDTH-1:229*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(3),
		.CELL_Z(3)
	)
	Pos_Cache_7_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[231*3*DATA_WIDTH-1:230*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(3),
		.CELL_Z(4)
	)
	Pos_Cache_7_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[232*3*DATA_WIDTH-1:231*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(3),
		.CELL_Z(5)
	)
	Pos_Cache_7_3_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[233*3*DATA_WIDTH-1:232*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(3),
		.CELL_Z(6)
	)
	Pos_Cache_7_3_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[234*3*DATA_WIDTH-1:233*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(4),
		.CELL_Z(1)
	)
	Pos_Cache_7_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[235*3*DATA_WIDTH-1:234*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(4),
		.CELL_Z(2)
	)
	Pos_Cache_7_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[236*3*DATA_WIDTH-1:235*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(4),
		.CELL_Z(3)
	)
	Pos_Cache_7_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[237*3*DATA_WIDTH-1:236*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(4),
		.CELL_Z(4)
	)
	Pos_Cache_7_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[238*3*DATA_WIDTH-1:237*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(4),
		.CELL_Z(5)
	)
	Pos_Cache_7_4_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[239*3*DATA_WIDTH-1:238*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(4),
		.CELL_Z(6)
	)
	Pos_Cache_7_4_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[240*3*DATA_WIDTH-1:239*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(5),
		.CELL_Z(1)
	)
	Pos_Cache_7_5_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[241*3*DATA_WIDTH-1:240*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(5),
		.CELL_Z(2)
	)
	Pos_Cache_7_5_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[242*3*DATA_WIDTH-1:241*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(5),
		.CELL_Z(3)
	)
	Pos_Cache_7_5_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[243*3*DATA_WIDTH-1:242*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(5),
		.CELL_Z(4)
	)
	Pos_Cache_7_5_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[244*3*DATA_WIDTH-1:243*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(5),
		.CELL_Z(5)
	)
	Pos_Cache_7_5_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[245*3*DATA_WIDTH-1:244*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(5),
		.CELL_Z(6)
	)
	Pos_Cache_7_5_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[246*3*DATA_WIDTH-1:245*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(6),
		.CELL_Z(1)
	)
	Pos_Cache_7_6_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[247*3*DATA_WIDTH-1:246*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(6),
		.CELL_Z(2)
	)
	Pos_Cache_7_6_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[248*3*DATA_WIDTH-1:247*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(6),
		.CELL_Z(3)
	)
	Pos_Cache_7_6_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[249*3*DATA_WIDTH-1:248*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(6),
		.CELL_Z(4)
	)
	Pos_Cache_7_6_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[250*3*DATA_WIDTH-1:249*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(6),
		.CELL_Z(5)
	)
	Pos_Cache_7_6_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[251*3*DATA_WIDTH-1:250*3*DATA_WIDTH])
	);

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(6),
		.CELL_Z(6)
	)
	Pos_Cache_7_6_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),								// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),									// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[252*3*DATA_WIDTH-1:251*3*DATA_WIDTH])
	);

	///////////////////////////////////////////////////////////////////////////////////////////////
	// Force cache
	// Each cell has an independent cache, MSB -> LSB:{Force_Z, Force_Y, Force_X}
	// The force Serve as the buffer to hold evaluated force values during evaluation
	// The initial force value is 0
	// When new force value arrives, it will accumulate to the current stored value
	///////////////////////////////////////////////////////////////////////////////////////////////
	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_1_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[0]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[1*PARTICLE_ID_WIDTH-1:0*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[0])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_1_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[1]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[2*PARTICLE_ID_WIDTH-1:1*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[1])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_1_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[2]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[3*PARTICLE_ID_WIDTH-1:2*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[2])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_1_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[3]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[4*PARTICLE_ID_WIDTH-1:3*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[3])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_1_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[4]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[5*PARTICLE_ID_WIDTH-1:4*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[4])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_1_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[5]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[6*PARTICLE_ID_WIDTH-1:5*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[5])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_2_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[6]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[7*PARTICLE_ID_WIDTH-1:6*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[6])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_2_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[7]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[8*PARTICLE_ID_WIDTH-1:7*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[7])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_2_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[8]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[9*3*DATA_WIDTH-1:8*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[9*PARTICLE_ID_WIDTH-1:8*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[8])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_2_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[9]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[10*3*DATA_WIDTH-1:9*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[10*PARTICLE_ID_WIDTH-1:9*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[9])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_2_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[10]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[11*3*DATA_WIDTH-1:10*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[11*PARTICLE_ID_WIDTH-1:10*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[10])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_2_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[11]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[12*3*DATA_WIDTH-1:11*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[12*PARTICLE_ID_WIDTH-1:11*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[11])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_3_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[12]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[13*3*DATA_WIDTH-1:12*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[13*PARTICLE_ID_WIDTH-1:12*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[12])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_3_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[13]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[14*3*DATA_WIDTH-1:13*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[14*PARTICLE_ID_WIDTH-1:13*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[13])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_3_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[14]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[15*3*DATA_WIDTH-1:14*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[15*PARTICLE_ID_WIDTH-1:14*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[14])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_3_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[15]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[16*3*DATA_WIDTH-1:15*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[16*PARTICLE_ID_WIDTH-1:15*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[15])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_3_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[16]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[17*PARTICLE_ID_WIDTH-1:16*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[16])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_3_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[17]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[18*PARTICLE_ID_WIDTH-1:17*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[17])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_4_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[18]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[19*PARTICLE_ID_WIDTH-1:18*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[18])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_4_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[19]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[20*PARTICLE_ID_WIDTH-1:19*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[19])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_4_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[20]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[21*PARTICLE_ID_WIDTH-1:20*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[20])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_4_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[21]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[22*PARTICLE_ID_WIDTH-1:21*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[21])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_4_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[22]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[23*PARTICLE_ID_WIDTH-1:22*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[22])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_4_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[23]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[24*PARTICLE_ID_WIDTH-1:23*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[23])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(5),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_5_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[24]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[25*3*DATA_WIDTH-1:24*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[25*PARTICLE_ID_WIDTH-1:24*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[24])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(5),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_5_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[25]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[26*3*DATA_WIDTH-1:25*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[26*PARTICLE_ID_WIDTH-1:25*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[25])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(5),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_5_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[26]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[27*3*DATA_WIDTH-1:26*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[27*PARTICLE_ID_WIDTH-1:26*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[26])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(5),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_5_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[27]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[28*3*DATA_WIDTH-1:27*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[28*PARTICLE_ID_WIDTH-1:27*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[27])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(5),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_5_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[28]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[29*PARTICLE_ID_WIDTH-1:28*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[28])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(5),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_5_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[29]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[30*PARTICLE_ID_WIDTH-1:29*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[29])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(6),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_6_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[30]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[31*PARTICLE_ID_WIDTH-1:30*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[30])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(6),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_6_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[31]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[32*PARTICLE_ID_WIDTH-1:31*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[31])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(6),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_6_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[32]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[33*3*DATA_WIDTH-1:32*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[33*PARTICLE_ID_WIDTH-1:32*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[32])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(6),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_6_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[33]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[34*3*DATA_WIDTH-1:33*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[34*PARTICLE_ID_WIDTH-1:33*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[33])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(6),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_6_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[34]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[35*3*DATA_WIDTH-1:34*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[35*PARTICLE_ID_WIDTH-1:34*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[34])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(1),
		.CELL_Y(6),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_1_6_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[35]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[36*3*DATA_WIDTH-1:35*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[36*PARTICLE_ID_WIDTH-1:35*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[35])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_1_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[36]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[37*3*DATA_WIDTH-1:36*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[37*PARTICLE_ID_WIDTH-1:36*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[36])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_1_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[37]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[38*3*DATA_WIDTH-1:37*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[38*PARTICLE_ID_WIDTH-1:37*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[37])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_1_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[38]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[39*3*DATA_WIDTH-1:38*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[39*PARTICLE_ID_WIDTH-1:38*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[38])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_1_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[39]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[40*3*DATA_WIDTH-1:39*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[40*PARTICLE_ID_WIDTH-1:39*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[39])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_1_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[40]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[41*3*DATA_WIDTH-1:40*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[41*PARTICLE_ID_WIDTH-1:40*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[40])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_1_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[41]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[42*3*DATA_WIDTH-1:41*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[42*PARTICLE_ID_WIDTH-1:41*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[41])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_2_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[42]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[43*3*DATA_WIDTH-1:42*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[43*PARTICLE_ID_WIDTH-1:42*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[42])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_2_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[43]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[44*3*DATA_WIDTH-1:43*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[44*PARTICLE_ID_WIDTH-1:43*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[43])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_2_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[44]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[45*3*DATA_WIDTH-1:44*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[45*PARTICLE_ID_WIDTH-1:44*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[44])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_2_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[45]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[46*3*DATA_WIDTH-1:45*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[46*PARTICLE_ID_WIDTH-1:45*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[45])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_2_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[46]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[47*3*DATA_WIDTH-1:46*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[47*PARTICLE_ID_WIDTH-1:46*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[46])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_2_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[47]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[48*3*DATA_WIDTH-1:47*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[48*PARTICLE_ID_WIDTH-1:47*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[47])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_3_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[48]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[49*3*DATA_WIDTH-1:48*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[49*PARTICLE_ID_WIDTH-1:48*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[48])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_3_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[49]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[50*3*DATA_WIDTH-1:49*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[50*PARTICLE_ID_WIDTH-1:49*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[49])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_3_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[50]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[51*3*DATA_WIDTH-1:50*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[51*PARTICLE_ID_WIDTH-1:50*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[50])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_3_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[51]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[52*3*DATA_WIDTH-1:51*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[52*PARTICLE_ID_WIDTH-1:51*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[51])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_3_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[52]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[53*3*DATA_WIDTH-1:52*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[53*PARTICLE_ID_WIDTH-1:52*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[52])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_3_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[53]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[54*3*DATA_WIDTH-1:53*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[54*PARTICLE_ID_WIDTH-1:53*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[53])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_4_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[54]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[55*3*DATA_WIDTH-1:54*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[55*PARTICLE_ID_WIDTH-1:54*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[54])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_4_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[55]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[56*3*DATA_WIDTH-1:55*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[56*PARTICLE_ID_WIDTH-1:55*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[55])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_4_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[56]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[57*3*DATA_WIDTH-1:56*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[57*PARTICLE_ID_WIDTH-1:56*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[56])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_4_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[57]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[58*3*DATA_WIDTH-1:57*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[58*PARTICLE_ID_WIDTH-1:57*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[57])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_4_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[58]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[59*3*DATA_WIDTH-1:58*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[59*PARTICLE_ID_WIDTH-1:58*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[58])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_4_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[59]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[60*3*DATA_WIDTH-1:59*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[60*PARTICLE_ID_WIDTH-1:59*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[59])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(5),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_5_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[60]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[61*3*DATA_WIDTH-1:60*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[61*PARTICLE_ID_WIDTH-1:60*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[60])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(5),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_5_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[61]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[62*3*DATA_WIDTH-1:61*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[62*PARTICLE_ID_WIDTH-1:61*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[61])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(5),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_5_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[62]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[63*3*DATA_WIDTH-1:62*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[63*PARTICLE_ID_WIDTH-1:62*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[62])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(5),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_5_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[63]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[64*3*DATA_WIDTH-1:63*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[64*PARTICLE_ID_WIDTH-1:63*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[63])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(5),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_5_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[64]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[65*3*DATA_WIDTH-1:64*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[65*PARTICLE_ID_WIDTH-1:64*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[64])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(5),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_5_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[65]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[66*3*DATA_WIDTH-1:65*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[66*PARTICLE_ID_WIDTH-1:65*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[65])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(6),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_6_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[66]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[67*3*DATA_WIDTH-1:66*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[67*PARTICLE_ID_WIDTH-1:66*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[66])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(6),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_6_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[67]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[68*3*DATA_WIDTH-1:67*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[68*PARTICLE_ID_WIDTH-1:67*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[67])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(6),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_6_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[68]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[69*3*DATA_WIDTH-1:68*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[69*PARTICLE_ID_WIDTH-1:68*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[68])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(6),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_6_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[69]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[70*3*DATA_WIDTH-1:69*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[70*PARTICLE_ID_WIDTH-1:69*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[69])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(6),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_6_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[70]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[71*3*DATA_WIDTH-1:70*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[71*PARTICLE_ID_WIDTH-1:70*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[70])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(2),
		.CELL_Y(6),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_2_6_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[71]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[72*3*DATA_WIDTH-1:71*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[72*PARTICLE_ID_WIDTH-1:71*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[71])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_1_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[72]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[73*3*DATA_WIDTH-1:72*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[73*PARTICLE_ID_WIDTH-1:72*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[72])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_1_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[73]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[74*3*DATA_WIDTH-1:73*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[74*PARTICLE_ID_WIDTH-1:73*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[73])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_1_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[74]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[75*3*DATA_WIDTH-1:74*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[75*PARTICLE_ID_WIDTH-1:74*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[74])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_1_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[75]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[76*3*DATA_WIDTH-1:75*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[76*PARTICLE_ID_WIDTH-1:75*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[75])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_1_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[76]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[77*3*DATA_WIDTH-1:76*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[77*PARTICLE_ID_WIDTH-1:76*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[76])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_1_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[77]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[78*3*DATA_WIDTH-1:77*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[78*PARTICLE_ID_WIDTH-1:77*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[77])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_2_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[78]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[79*3*DATA_WIDTH-1:78*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[79*PARTICLE_ID_WIDTH-1:78*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[78])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_2_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[79]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[80*3*DATA_WIDTH-1:79*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[80*PARTICLE_ID_WIDTH-1:79*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[79])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_2_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[80]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[81*3*DATA_WIDTH-1:80*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[81*PARTICLE_ID_WIDTH-1:80*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[80])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_2_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[81]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[82*3*DATA_WIDTH-1:81*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[82*PARTICLE_ID_WIDTH-1:81*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[81])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_2_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[82]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[83*3*DATA_WIDTH-1:82*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[83*PARTICLE_ID_WIDTH-1:82*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[82])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_2_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[83]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[84*3*DATA_WIDTH-1:83*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[84*PARTICLE_ID_WIDTH-1:83*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[83])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_3_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[84]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[85*3*DATA_WIDTH-1:84*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[85*PARTICLE_ID_WIDTH-1:84*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[84])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_3_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[85]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[86*3*DATA_WIDTH-1:85*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[86*PARTICLE_ID_WIDTH-1:85*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[85])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_3_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[86]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[87*3*DATA_WIDTH-1:86*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[87*PARTICLE_ID_WIDTH-1:86*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[86])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_3_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[87]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[88*3*DATA_WIDTH-1:87*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[88*PARTICLE_ID_WIDTH-1:87*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[87])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_3_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[88]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[89*3*DATA_WIDTH-1:88*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[89*PARTICLE_ID_WIDTH-1:88*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[88])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_3_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[89]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[90*3*DATA_WIDTH-1:89*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[90*PARTICLE_ID_WIDTH-1:89*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[89])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_4_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[90]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[91*3*DATA_WIDTH-1:90*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[91*PARTICLE_ID_WIDTH-1:90*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[90])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_4_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[91]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[92*3*DATA_WIDTH-1:91*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[92*PARTICLE_ID_WIDTH-1:91*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[91])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_4_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[92]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[93*3*DATA_WIDTH-1:92*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[93*PARTICLE_ID_WIDTH-1:92*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[92])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_4_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[93]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[94*3*DATA_WIDTH-1:93*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[94*PARTICLE_ID_WIDTH-1:93*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[93])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_4_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[94]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[95*3*DATA_WIDTH-1:94*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[95*PARTICLE_ID_WIDTH-1:94*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[94])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_4_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[95]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[96*3*DATA_WIDTH-1:95*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[96*PARTICLE_ID_WIDTH-1:95*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[95])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(5),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_5_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[96]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[97*3*DATA_WIDTH-1:96*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[97*PARTICLE_ID_WIDTH-1:96*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[96])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(5),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_5_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[97]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[98*3*DATA_WIDTH-1:97*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[98*PARTICLE_ID_WIDTH-1:97*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[97])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(5),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_5_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[98]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[99*3*DATA_WIDTH-1:98*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[99*PARTICLE_ID_WIDTH-1:98*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[98])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(5),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_5_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[99]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[100*3*DATA_WIDTH-1:99*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[100*PARTICLE_ID_WIDTH-1:99*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[99])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(5),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_5_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[100]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[101*3*DATA_WIDTH-1:100*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[101*PARTICLE_ID_WIDTH-1:100*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[100])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(5),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_5_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[101]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[102*3*DATA_WIDTH-1:101*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[102*PARTICLE_ID_WIDTH-1:101*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[101])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(6),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_6_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[102]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[103*3*DATA_WIDTH-1:102*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[103*PARTICLE_ID_WIDTH-1:102*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[102])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(6),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_6_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[103]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[104*3*DATA_WIDTH-1:103*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[104*PARTICLE_ID_WIDTH-1:103*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[103])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(6),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_6_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[104]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[105*3*DATA_WIDTH-1:104*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[105*PARTICLE_ID_WIDTH-1:104*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[104])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(6),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_6_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[105]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[106*3*DATA_WIDTH-1:105*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[106*PARTICLE_ID_WIDTH-1:105*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[105])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(6),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_6_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[106]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[107*3*DATA_WIDTH-1:106*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[107*PARTICLE_ID_WIDTH-1:106*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[106])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(3),
		.CELL_Y(6),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_3_6_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[107]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[108*3*DATA_WIDTH-1:107*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[108*PARTICLE_ID_WIDTH-1:107*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[107])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_1_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[108]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[109*3*DATA_WIDTH-1:108*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[109*PARTICLE_ID_WIDTH-1:108*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[108])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_1_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[109]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[110*3*DATA_WIDTH-1:109*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[110*PARTICLE_ID_WIDTH-1:109*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[109])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_1_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[110]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[111*3*DATA_WIDTH-1:110*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[111*PARTICLE_ID_WIDTH-1:110*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[110])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_1_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[111]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[112*3*DATA_WIDTH-1:111*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[112*PARTICLE_ID_WIDTH-1:111*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[111])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_1_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[112]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[113*3*DATA_WIDTH-1:112*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[113*PARTICLE_ID_WIDTH-1:112*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[112])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_1_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[113]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[114*3*DATA_WIDTH-1:113*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[114*PARTICLE_ID_WIDTH-1:113*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[113])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_2_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[114]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[115*3*DATA_WIDTH-1:114*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[115*PARTICLE_ID_WIDTH-1:114*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[114])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_2_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[115]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[116*3*DATA_WIDTH-1:115*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[116*PARTICLE_ID_WIDTH-1:115*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[115])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_2_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[116]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[117*3*DATA_WIDTH-1:116*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[117*PARTICLE_ID_WIDTH-1:116*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[116])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_2_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[117]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[118*3*DATA_WIDTH-1:117*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[118*PARTICLE_ID_WIDTH-1:117*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[117])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_2_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[118]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[119*3*DATA_WIDTH-1:118*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[119*PARTICLE_ID_WIDTH-1:118*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[118])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_2_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[119]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[120*3*DATA_WIDTH-1:119*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[120*PARTICLE_ID_WIDTH-1:119*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[119])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_3_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[120]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[121*3*DATA_WIDTH-1:120*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[121*PARTICLE_ID_WIDTH-1:120*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[120])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_3_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[121]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[122*3*DATA_WIDTH-1:121*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[122*PARTICLE_ID_WIDTH-1:121*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[121])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_3_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[122]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[123*3*DATA_WIDTH-1:122*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[123*PARTICLE_ID_WIDTH-1:122*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[122])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_3_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[123]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[124*3*DATA_WIDTH-1:123*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[124*PARTICLE_ID_WIDTH-1:123*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[123])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_3_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[124]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[125*3*DATA_WIDTH-1:124*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[125*PARTICLE_ID_WIDTH-1:124*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[124])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_3_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[125]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[126*3*DATA_WIDTH-1:125*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[126*PARTICLE_ID_WIDTH-1:125*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[125])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_4_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[126]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[127*3*DATA_WIDTH-1:126*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[127*PARTICLE_ID_WIDTH-1:126*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[126])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_4_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[127]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[128*3*DATA_WIDTH-1:127*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[128*PARTICLE_ID_WIDTH-1:127*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[127])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_4_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[128]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[129*3*DATA_WIDTH-1:128*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[129*PARTICLE_ID_WIDTH-1:128*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[128])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_4_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[129]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[130*3*DATA_WIDTH-1:129*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[130*PARTICLE_ID_WIDTH-1:129*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[129])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_4_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[130]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[131*3*DATA_WIDTH-1:130*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[131*PARTICLE_ID_WIDTH-1:130*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[130])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_4_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[131]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[132*3*DATA_WIDTH-1:131*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[132*PARTICLE_ID_WIDTH-1:131*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[131])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(5),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_5_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[132]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[133*3*DATA_WIDTH-1:132*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[133*PARTICLE_ID_WIDTH-1:132*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[132])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(5),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_5_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[133]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[134*3*DATA_WIDTH-1:133*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[134*PARTICLE_ID_WIDTH-1:133*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[133])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(5),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_5_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[134]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[135*3*DATA_WIDTH-1:134*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[135*PARTICLE_ID_WIDTH-1:134*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[134])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(5),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_5_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[135]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[136*3*DATA_WIDTH-1:135*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[136*PARTICLE_ID_WIDTH-1:135*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[135])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(5),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_5_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[136]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[137*3*DATA_WIDTH-1:136*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[137*PARTICLE_ID_WIDTH-1:136*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[136])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(5),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_5_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[137]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[138*3*DATA_WIDTH-1:137*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[138*PARTICLE_ID_WIDTH-1:137*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[137])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(6),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_6_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[138]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[139*3*DATA_WIDTH-1:138*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[139*PARTICLE_ID_WIDTH-1:138*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[138])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(6),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_6_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[139]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[140*3*DATA_WIDTH-1:139*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[140*PARTICLE_ID_WIDTH-1:139*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[139])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(6),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_6_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[140]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[141*3*DATA_WIDTH-1:140*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[141*PARTICLE_ID_WIDTH-1:140*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[140])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(6),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_6_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[141]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[142*3*DATA_WIDTH-1:141*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[142*PARTICLE_ID_WIDTH-1:141*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[141])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(6),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_6_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[142]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[143*3*DATA_WIDTH-1:142*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[143*PARTICLE_ID_WIDTH-1:142*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[142])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(4),
		.CELL_Y(6),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_4_6_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[143]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[144*3*DATA_WIDTH-1:143*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[144*PARTICLE_ID_WIDTH-1:143*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[143])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(1),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_1_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[144]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[145*3*DATA_WIDTH-1:144*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[145*PARTICLE_ID_WIDTH-1:144*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[144])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(1),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_1_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[145]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[146*3*DATA_WIDTH-1:145*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[146*PARTICLE_ID_WIDTH-1:145*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[145])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(1),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_1_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[146]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[147*3*DATA_WIDTH-1:146*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[147*PARTICLE_ID_WIDTH-1:146*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[146])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(1),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_1_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[147]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[148*3*DATA_WIDTH-1:147*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[148*PARTICLE_ID_WIDTH-1:147*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[147])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(1),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_1_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[148]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[149*3*DATA_WIDTH-1:148*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[149*PARTICLE_ID_WIDTH-1:148*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[148])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(1),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_1_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[149]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[150*3*DATA_WIDTH-1:149*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[150*PARTICLE_ID_WIDTH-1:149*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[149])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(2),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_2_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[150]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[151*3*DATA_WIDTH-1:150*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[151*PARTICLE_ID_WIDTH-1:150*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[150])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(2),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_2_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[151]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[152*3*DATA_WIDTH-1:151*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[152*PARTICLE_ID_WIDTH-1:151*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[151])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(2),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_2_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[152]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[153*3*DATA_WIDTH-1:152*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[153*PARTICLE_ID_WIDTH-1:152*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[152])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(2),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_2_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[153]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[154*3*DATA_WIDTH-1:153*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[154*PARTICLE_ID_WIDTH-1:153*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[153])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(2),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_2_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[154]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[155*3*DATA_WIDTH-1:154*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[155*PARTICLE_ID_WIDTH-1:154*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[154])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(2),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_2_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[155]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[156*3*DATA_WIDTH-1:155*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[156*PARTICLE_ID_WIDTH-1:155*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[155])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(3),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_3_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[156]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[157*3*DATA_WIDTH-1:156*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[157*PARTICLE_ID_WIDTH-1:156*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[156])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(3),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_3_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[157]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[158*3*DATA_WIDTH-1:157*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[158*PARTICLE_ID_WIDTH-1:157*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[157])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(3),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_3_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[158]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[159*3*DATA_WIDTH-1:158*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[159*PARTICLE_ID_WIDTH-1:158*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[158])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(3),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_3_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[159]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[160*3*DATA_WIDTH-1:159*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[160*PARTICLE_ID_WIDTH-1:159*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[159])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(3),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_3_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[160]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[161*3*DATA_WIDTH-1:160*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[161*PARTICLE_ID_WIDTH-1:160*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[160])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(3),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_3_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[161]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[162*3*DATA_WIDTH-1:161*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[162*PARTICLE_ID_WIDTH-1:161*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[161])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(4),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_4_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[162]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[163*3*DATA_WIDTH-1:162*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[163*PARTICLE_ID_WIDTH-1:162*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[162])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(4),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_4_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[163]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[164*3*DATA_WIDTH-1:163*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[164*PARTICLE_ID_WIDTH-1:163*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[163])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(4),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_4_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[164]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[165*3*DATA_WIDTH-1:164*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[165*PARTICLE_ID_WIDTH-1:164*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[164])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(4),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_4_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[165]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[166*3*DATA_WIDTH-1:165*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[166*PARTICLE_ID_WIDTH-1:165*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[165])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(4),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_4_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[166]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[167*3*DATA_WIDTH-1:166*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[167*PARTICLE_ID_WIDTH-1:166*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[166])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(4),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_4_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[167]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[168*3*DATA_WIDTH-1:167*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[168*PARTICLE_ID_WIDTH-1:167*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[167])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(5),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_5_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[168]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[169*3*DATA_WIDTH-1:168*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[169*PARTICLE_ID_WIDTH-1:168*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[168])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(5),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_5_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[169]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[170*3*DATA_WIDTH-1:169*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[170*PARTICLE_ID_WIDTH-1:169*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[169])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(5),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_5_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[170]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[171*3*DATA_WIDTH-1:170*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[171*PARTICLE_ID_WIDTH-1:170*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[170])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(5),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_5_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[171]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[172*3*DATA_WIDTH-1:171*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[172*PARTICLE_ID_WIDTH-1:171*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[171])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(5),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_5_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[172]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[173*3*DATA_WIDTH-1:172*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[173*PARTICLE_ID_WIDTH-1:172*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[172])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(5),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_5_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[173]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[174*3*DATA_WIDTH-1:173*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[174*PARTICLE_ID_WIDTH-1:173*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[173])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(6),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_6_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[174]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[175*3*DATA_WIDTH-1:174*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[175*PARTICLE_ID_WIDTH-1:174*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[174])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(6),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_6_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[175]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[176*3*DATA_WIDTH-1:175*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[176*PARTICLE_ID_WIDTH-1:175*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[175])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(6),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_6_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[176]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[177*3*DATA_WIDTH-1:176*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[177*PARTICLE_ID_WIDTH-1:176*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[176])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(6),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_6_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[177]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[178*3*DATA_WIDTH-1:177*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[178*PARTICLE_ID_WIDTH-1:177*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[177])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(6),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_6_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[178]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[179*3*DATA_WIDTH-1:178*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[179*PARTICLE_ID_WIDTH-1:178*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[178])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(5),
		.CELL_Y(6),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_5_6_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[179]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[180*3*DATA_WIDTH-1:179*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[180*PARTICLE_ID_WIDTH-1:179*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[179])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(1),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_1_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[180]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[181*3*DATA_WIDTH-1:180*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[181*PARTICLE_ID_WIDTH-1:180*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[180])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(1),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_1_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[181]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[182*3*DATA_WIDTH-1:181*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[182*PARTICLE_ID_WIDTH-1:181*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[181])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(1),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_1_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[182]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[183*3*DATA_WIDTH-1:182*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[183*PARTICLE_ID_WIDTH-1:182*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[182])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(1),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_1_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[183]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[184*3*DATA_WIDTH-1:183*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[184*PARTICLE_ID_WIDTH-1:183*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[183])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(1),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_1_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[184]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[185*3*DATA_WIDTH-1:184*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[185*PARTICLE_ID_WIDTH-1:184*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[184])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(1),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_1_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[185]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[186*3*DATA_WIDTH-1:185*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[186*PARTICLE_ID_WIDTH-1:185*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[185])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(2),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_2_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[186]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[187*3*DATA_WIDTH-1:186*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[187*PARTICLE_ID_WIDTH-1:186*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[186])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(2),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_2_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[187]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[188*3*DATA_WIDTH-1:187*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[188*PARTICLE_ID_WIDTH-1:187*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[187])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(2),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_2_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[188]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[189*3*DATA_WIDTH-1:188*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[189*PARTICLE_ID_WIDTH-1:188*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[188])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(2),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_2_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[189]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[190*3*DATA_WIDTH-1:189*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[190*PARTICLE_ID_WIDTH-1:189*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[189])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(2),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_2_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[190]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[191*3*DATA_WIDTH-1:190*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[191*PARTICLE_ID_WIDTH-1:190*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[190])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(2),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_2_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[191]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[192*3*DATA_WIDTH-1:191*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[192*PARTICLE_ID_WIDTH-1:191*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[191])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(3),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_3_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[192]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[193*3*DATA_WIDTH-1:192*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[193*PARTICLE_ID_WIDTH-1:192*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[192])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(3),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_3_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[193]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[194*3*DATA_WIDTH-1:193*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[194*PARTICLE_ID_WIDTH-1:193*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[193])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(3),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_3_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[194]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[195*3*DATA_WIDTH-1:194*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[195*PARTICLE_ID_WIDTH-1:194*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[194])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(3),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_3_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[195]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[196*3*DATA_WIDTH-1:195*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[196*PARTICLE_ID_WIDTH-1:195*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[195])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(3),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_3_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[196]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[197*3*DATA_WIDTH-1:196*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[197*PARTICLE_ID_WIDTH-1:196*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[196])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(3),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_3_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[197]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[198*3*DATA_WIDTH-1:197*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[198*PARTICLE_ID_WIDTH-1:197*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[197])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(4),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_4_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[198]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[199*3*DATA_WIDTH-1:198*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[199*PARTICLE_ID_WIDTH-1:198*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[198])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(4),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_4_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[199]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[200*3*DATA_WIDTH-1:199*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[200*PARTICLE_ID_WIDTH-1:199*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[199])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(4),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_4_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[200]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[201*3*DATA_WIDTH-1:200*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[201*PARTICLE_ID_WIDTH-1:200*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[200])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(4),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_4_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[201]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[202*3*DATA_WIDTH-1:201*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[202*PARTICLE_ID_WIDTH-1:201*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[201])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(4),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_4_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[202]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[203*3*DATA_WIDTH-1:202*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[203*PARTICLE_ID_WIDTH-1:202*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[202])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(4),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_4_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[203]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[204*3*DATA_WIDTH-1:203*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[204*PARTICLE_ID_WIDTH-1:203*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[203])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(5),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_5_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[204]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[205*3*DATA_WIDTH-1:204*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[205*PARTICLE_ID_WIDTH-1:204*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[204])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(5),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_5_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[205]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[206*3*DATA_WIDTH-1:205*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[206*PARTICLE_ID_WIDTH-1:205*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[205])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(5),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_5_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[206]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[207*3*DATA_WIDTH-1:206*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[207*PARTICLE_ID_WIDTH-1:206*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[206])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(5),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_5_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[207]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[208*3*DATA_WIDTH-1:207*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[208*PARTICLE_ID_WIDTH-1:207*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[207])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(5),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_5_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[208]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[209*3*DATA_WIDTH-1:208*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[209*PARTICLE_ID_WIDTH-1:208*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[208])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(5),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_5_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[209]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[210*3*DATA_WIDTH-1:209*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[210*PARTICLE_ID_WIDTH-1:209*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[209])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(6),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_6_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[210]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[211*3*DATA_WIDTH-1:210*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[211*PARTICLE_ID_WIDTH-1:210*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[210])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(6),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_6_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[211]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[212*3*DATA_WIDTH-1:211*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[212*PARTICLE_ID_WIDTH-1:211*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[211])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(6),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_6_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[212]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[213*3*DATA_WIDTH-1:212*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[213*PARTICLE_ID_WIDTH-1:212*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[212])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(6),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_6_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[213]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[214*3*DATA_WIDTH-1:213*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[214*PARTICLE_ID_WIDTH-1:213*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[213])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(6),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_6_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[214]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[215*3*DATA_WIDTH-1:214*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[215*PARTICLE_ID_WIDTH-1:214*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[214])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(6),
		.CELL_Y(6),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_6_6_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[215]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[216*3*DATA_WIDTH-1:215*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[216*PARTICLE_ID_WIDTH-1:215*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[215])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(1),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_1_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[216]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[217*3*DATA_WIDTH-1:216*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[217*PARTICLE_ID_WIDTH-1:216*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[216])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(1),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_1_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[217]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[218*3*DATA_WIDTH-1:217*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[218*PARTICLE_ID_WIDTH-1:217*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[217])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(1),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_1_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[218]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[219*3*DATA_WIDTH-1:218*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[219*PARTICLE_ID_WIDTH-1:218*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[218])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(1),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_1_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[219]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[220*3*DATA_WIDTH-1:219*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[220*PARTICLE_ID_WIDTH-1:219*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[219])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(1),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_1_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[220]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[221*3*DATA_WIDTH-1:220*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[221*PARTICLE_ID_WIDTH-1:220*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[220])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(1),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_1_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[221]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[222*3*DATA_WIDTH-1:221*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[222*PARTICLE_ID_WIDTH-1:221*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[221])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(2),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_2_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[222]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[223*3*DATA_WIDTH-1:222*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[223*PARTICLE_ID_WIDTH-1:222*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[222])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(2),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_2_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[223]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[224*3*DATA_WIDTH-1:223*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[224*PARTICLE_ID_WIDTH-1:223*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[223])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(2),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_2_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[224]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[225*3*DATA_WIDTH-1:224*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[225*PARTICLE_ID_WIDTH-1:224*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[224])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(2),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_2_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[225]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[226*3*DATA_WIDTH-1:225*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[226*PARTICLE_ID_WIDTH-1:225*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[225])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(2),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_2_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[226]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[227*3*DATA_WIDTH-1:226*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[227*PARTICLE_ID_WIDTH-1:226*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[226])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(2),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_2_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[227]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[228*3*DATA_WIDTH-1:227*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[228*PARTICLE_ID_WIDTH-1:227*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[227])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(3),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_3_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[228]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[229*3*DATA_WIDTH-1:228*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[229*PARTICLE_ID_WIDTH-1:228*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[228])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(3),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_3_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[229]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[230*3*DATA_WIDTH-1:229*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[230*PARTICLE_ID_WIDTH-1:229*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[229])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(3),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_3_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[230]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[231*3*DATA_WIDTH-1:230*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[231*PARTICLE_ID_WIDTH-1:230*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[230])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(3),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_3_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[231]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[232*3*DATA_WIDTH-1:231*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[232*PARTICLE_ID_WIDTH-1:231*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[231])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(3),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_3_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[232]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[233*3*DATA_WIDTH-1:232*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[233*PARTICLE_ID_WIDTH-1:232*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[232])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(3),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_3_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[233]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[234*3*DATA_WIDTH-1:233*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[234*PARTICLE_ID_WIDTH-1:233*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[233])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(4),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_4_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[234]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[235*3*DATA_WIDTH-1:234*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[235*PARTICLE_ID_WIDTH-1:234*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[234])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(4),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_4_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[235]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[236*3*DATA_WIDTH-1:235*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[236*PARTICLE_ID_WIDTH-1:235*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[235])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(4),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_4_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[236]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[237*3*DATA_WIDTH-1:236*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[237*PARTICLE_ID_WIDTH-1:236*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[236])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(4),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_4_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[237]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[238*3*DATA_WIDTH-1:237*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[238*PARTICLE_ID_WIDTH-1:237*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[237])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(4),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_4_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[238]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[239*3*DATA_WIDTH-1:238*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[239*PARTICLE_ID_WIDTH-1:238*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[238])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(4),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_4_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[239]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[240*3*DATA_WIDTH-1:239*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[240*PARTICLE_ID_WIDTH-1:239*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[239])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(5),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_5_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[240]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[241*3*DATA_WIDTH-1:240*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[241*PARTICLE_ID_WIDTH-1:240*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[240])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(5),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_5_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[241]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[242*3*DATA_WIDTH-1:241*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[242*PARTICLE_ID_WIDTH-1:241*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[241])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(5),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_5_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[242]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[243*3*DATA_WIDTH-1:242*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[243*PARTICLE_ID_WIDTH-1:242*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[242])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(5),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_5_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[243]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[244*3*DATA_WIDTH-1:243*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[244*PARTICLE_ID_WIDTH-1:243*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[243])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(5),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_5_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[244]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[245*3*DATA_WIDTH-1:244*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[245*PARTICLE_ID_WIDTH-1:244*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[244])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(5),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_5_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[245]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[246*3*DATA_WIDTH-1:245*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[246*PARTICLE_ID_WIDTH-1:245*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[245])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(6),
		.CELL_Z(1),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_6_1
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[246]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[247*3*DATA_WIDTH-1:246*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[247*PARTICLE_ID_WIDTH-1:246*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[246])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(6),
		.CELL_Z(2),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_6_2
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[247]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[248*3*DATA_WIDTH-1:247*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[248*PARTICLE_ID_WIDTH-1:247*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[247])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(6),
		.CELL_Z(3),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_6_3
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[248]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[249*3*DATA_WIDTH-1:248*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[249*PARTICLE_ID_WIDTH-1:248*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[248])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(6),
		.CELL_Z(4),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_6_4
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[249]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[250*3*DATA_WIDTH-1:249*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[250*PARTICLE_ID_WIDTH-1:249*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[249])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(6),
		.CELL_Z(5),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_6_5
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[250]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[251*3*DATA_WIDTH-1:250*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[251*PARTICLE_ID_WIDTH-1:250*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[250])
	);

	Force_Write_Back_Controller
	#(
		.DATA_WIDTH(DATA_WIDTH),							// Data width of a single force value, 32-bit
		// Cell id this unit related to
		.CELL_X(7),
		.CELL_Y(6),
		.CELL_Z(6),
		// Force cache input buffer
		.FORCE_CACHE_BUFFER_DEPTH(FORCE_CACHE_BUFFER_DEPTH),
		.FORCE_CACHE_BUFFER_ADDR_WIDTH(FORCE_CACHE_BUFFER_ADDR_WIDTH),	// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
		// Dataset defined parameters
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.MAX_CELL_PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),		// The maximum # of particles can be in a cell
		.CELL_ADDR_WIDTH(CELL_ADDR_WIDTH),					// log(MAX_CELL_PARTICLE_NUM)
		.PARTICLE_ID_WIDTH(PARTICLE_ID_WIDTH)				// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
		
	)
	Force_Cache_7_6_6
	(
		.clk(clk),
		.rst(rst),
		// Cache input force
		.in_partial_force_valid(ref_forceoutput_valid),
		.in_particle_id(ref_particle_id),
		.in_partial_force({ref_LJ_Force_Z, ref_LJ_Force_Y, ref_LJ_Force_X}),
		// Cache output force
		.in_read_data_request(wire_motion_update_to_cache_read_force_request[251]),
		.in_cache_read_address(Motion_Update_force_read_addr),
		.out_partial_force(wire_cache_to_motion_update_partial_force[252*3*DATA_WIDTH-1:251*3*DATA_WIDTH]),
		.out_particle_id(wire_cache_to_motion_update_particle_id[252*PARTICLE_ID_WIDTH-1:251*PARTICLE_ID_WIDTH]),
		.out_cache_readout_valid(wire_cache_to_motion_update_partial_force_valid[251])
	);

	///////////////////////////////////////////////////////////////////////////////////////////////
	// Velocity cache
	// Each cell has an independent cache, MSB -> LSB:{vz, vy, vx}
	// The velocity cache provide the spped information for motion update units
	// The inital velocity information is initialized by a initilization file generated from scripts
	// Double buffer mechanism is implemented
	// During motion update process, the new evaluated speed information will write into the alternative cache
	// The read and write address and particle number information should be the same as the Position Cache
	///////////////////////////////////////////////////////////////////////////////////////////////
	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(1)
	)
	Velocity_Cache_1_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(2)
	)
	Velocity_Cache_1_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(3)
	)
	Velocity_Cache_1_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(4)
	)
	Velocity_Cache_1_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(5)
	)
	Velocity_Cache_1_1_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(6)
	)
	Velocity_Cache_1_1_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(1)
	)
	Velocity_Cache_1_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(2)
	)
	Velocity_Cache_1_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(3)
	)
	Velocity_Cache_1_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[9*3*DATA_WIDTH-1:8*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(4)
	)
	Velocity_Cache_1_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[10*3*DATA_WIDTH-1:9*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(5)
	)
	Velocity_Cache_1_2_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[11*3*DATA_WIDTH-1:10*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(6)
	)
	Velocity_Cache_1_2_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[12*3*DATA_WIDTH-1:11*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(1)
	)
	Velocity_Cache_1_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[13*3*DATA_WIDTH-1:12*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(2)
	)
	Velocity_Cache_1_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[14*3*DATA_WIDTH-1:13*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(3)
	)
	Velocity_Cache_1_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[15*3*DATA_WIDTH-1:14*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(4)
	)
	Velocity_Cache_1_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[16*3*DATA_WIDTH-1:15*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(5)
	)
	Velocity_Cache_1_3_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(6)
	)
	Velocity_Cache_1_3_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(1)
	)
	Velocity_Cache_1_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(2)
	)
	Velocity_Cache_1_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(3)
	)
	Velocity_Cache_1_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(4)
	)
	Velocity_Cache_1_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(5)
	)
	Velocity_Cache_1_4_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(6)
	)
	Velocity_Cache_1_4_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(5),
		.CELL_Z(1)
	)
	Velocity_Cache_1_5_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[25*3*DATA_WIDTH-1:24*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(5),
		.CELL_Z(2)
	)
	Velocity_Cache_1_5_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[26*3*DATA_WIDTH-1:25*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(5),
		.CELL_Z(3)
	)
	Velocity_Cache_1_5_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[27*3*DATA_WIDTH-1:26*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(5),
		.CELL_Z(4)
	)
	Velocity_Cache_1_5_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[28*3*DATA_WIDTH-1:27*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(5),
		.CELL_Z(5)
	)
	Velocity_Cache_1_5_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(5),
		.CELL_Z(6)
	)
	Velocity_Cache_1_5_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(6),
		.CELL_Z(1)
	)
	Velocity_Cache_1_6_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(6),
		.CELL_Z(2)
	)
	Velocity_Cache_1_6_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(6),
		.CELL_Z(3)
	)
	Velocity_Cache_1_6_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[33*3*DATA_WIDTH-1:32*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(6),
		.CELL_Z(4)
	)
	Velocity_Cache_1_6_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[34*3*DATA_WIDTH-1:33*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(6),
		.CELL_Z(5)
	)
	Velocity_Cache_1_6_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[35*3*DATA_WIDTH-1:34*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(6),
		.CELL_Z(6)
	)
	Velocity_Cache_1_6_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[36*3*DATA_WIDTH-1:35*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(1)
	)
	Velocity_Cache_2_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[37*3*DATA_WIDTH-1:36*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(2)
	)
	Velocity_Cache_2_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[38*3*DATA_WIDTH-1:37*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(3)
	)
	Velocity_Cache_2_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[39*3*DATA_WIDTH-1:38*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(4)
	)
	Velocity_Cache_2_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[40*3*DATA_WIDTH-1:39*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(5)
	)
	Velocity_Cache_2_1_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[41*3*DATA_WIDTH-1:40*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(6)
	)
	Velocity_Cache_2_1_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[42*3*DATA_WIDTH-1:41*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(1)
	)
	Velocity_Cache_2_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[43*3*DATA_WIDTH-1:42*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(2)
	)
	Velocity_Cache_2_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[44*3*DATA_WIDTH-1:43*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(3)
	)
	Velocity_Cache_2_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[45*3*DATA_WIDTH-1:44*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(4)
	)
	Velocity_Cache_2_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[46*3*DATA_WIDTH-1:45*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(5)
	)
	Velocity_Cache_2_2_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[47*3*DATA_WIDTH-1:46*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(6)
	)
	Velocity_Cache_2_2_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[48*3*DATA_WIDTH-1:47*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(1)
	)
	Velocity_Cache_2_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[49*3*DATA_WIDTH-1:48*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(2)
	)
	Velocity_Cache_2_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[50*3*DATA_WIDTH-1:49*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(3)
	)
	Velocity_Cache_2_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[51*3*DATA_WIDTH-1:50*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(4)
	)
	Velocity_Cache_2_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[52*3*DATA_WIDTH-1:51*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(5)
	)
	Velocity_Cache_2_3_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[53*3*DATA_WIDTH-1:52*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(6)
	)
	Velocity_Cache_2_3_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[54*3*DATA_WIDTH-1:53*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(1)
	)
	Velocity_Cache_2_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[55*3*DATA_WIDTH-1:54*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(2)
	)
	Velocity_Cache_2_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[56*3*DATA_WIDTH-1:55*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(3)
	)
	Velocity_Cache_2_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[57*3*DATA_WIDTH-1:56*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(4)
	)
	Velocity_Cache_2_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[58*3*DATA_WIDTH-1:57*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(5)
	)
	Velocity_Cache_2_4_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[59*3*DATA_WIDTH-1:58*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(6)
	)
	Velocity_Cache_2_4_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[60*3*DATA_WIDTH-1:59*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(5),
		.CELL_Z(1)
	)
	Velocity_Cache_2_5_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[61*3*DATA_WIDTH-1:60*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(5),
		.CELL_Z(2)
	)
	Velocity_Cache_2_5_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[62*3*DATA_WIDTH-1:61*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(5),
		.CELL_Z(3)
	)
	Velocity_Cache_2_5_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[63*3*DATA_WIDTH-1:62*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(5),
		.CELL_Z(4)
	)
	Velocity_Cache_2_5_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[64*3*DATA_WIDTH-1:63*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(5),
		.CELL_Z(5)
	)
	Velocity_Cache_2_5_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[65*3*DATA_WIDTH-1:64*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(5),
		.CELL_Z(6)
	)
	Velocity_Cache_2_5_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[66*3*DATA_WIDTH-1:65*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(6),
		.CELL_Z(1)
	)
	Velocity_Cache_2_6_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[67*3*DATA_WIDTH-1:66*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(6),
		.CELL_Z(2)
	)
	Velocity_Cache_2_6_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[68*3*DATA_WIDTH-1:67*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(6),
		.CELL_Z(3)
	)
	Velocity_Cache_2_6_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[69*3*DATA_WIDTH-1:68*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(6),
		.CELL_Z(4)
	)
	Velocity_Cache_2_6_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[70*3*DATA_WIDTH-1:69*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(6),
		.CELL_Z(5)
	)
	Velocity_Cache_2_6_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[71*3*DATA_WIDTH-1:70*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(6),
		.CELL_Z(6)
	)
	Velocity_Cache_2_6_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[72*3*DATA_WIDTH-1:71*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(1)
	)
	Velocity_Cache_3_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[73*3*DATA_WIDTH-1:72*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(2)
	)
	Velocity_Cache_3_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[74*3*DATA_WIDTH-1:73*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(3)
	)
	Velocity_Cache_3_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[75*3*DATA_WIDTH-1:74*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(4)
	)
	Velocity_Cache_3_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[76*3*DATA_WIDTH-1:75*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(5)
	)
	Velocity_Cache_3_1_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[77*3*DATA_WIDTH-1:76*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(6)
	)
	Velocity_Cache_3_1_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[78*3*DATA_WIDTH-1:77*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(1)
	)
	Velocity_Cache_3_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[79*3*DATA_WIDTH-1:78*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(2)
	)
	Velocity_Cache_3_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[80*3*DATA_WIDTH-1:79*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(3)
	)
	Velocity_Cache_3_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[81*3*DATA_WIDTH-1:80*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(4)
	)
	Velocity_Cache_3_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[82*3*DATA_WIDTH-1:81*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(5)
	)
	Velocity_Cache_3_2_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[83*3*DATA_WIDTH-1:82*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(6)
	)
	Velocity_Cache_3_2_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[84*3*DATA_WIDTH-1:83*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(1)
	)
	Velocity_Cache_3_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[85*3*DATA_WIDTH-1:84*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(2)
	)
	Velocity_Cache_3_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[86*3*DATA_WIDTH-1:85*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(3)
	)
	Velocity_Cache_3_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[87*3*DATA_WIDTH-1:86*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(4)
	)
	Velocity_Cache_3_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[88*3*DATA_WIDTH-1:87*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(5)
	)
	Velocity_Cache_3_3_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[89*3*DATA_WIDTH-1:88*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(6)
	)
	Velocity_Cache_3_3_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[90*3*DATA_WIDTH-1:89*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(1)
	)
	Velocity_Cache_3_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[91*3*DATA_WIDTH-1:90*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(2)
	)
	Velocity_Cache_3_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[92*3*DATA_WIDTH-1:91*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(3)
	)
	Velocity_Cache_3_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[93*3*DATA_WIDTH-1:92*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(4)
	)
	Velocity_Cache_3_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[94*3*DATA_WIDTH-1:93*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(5)
	)
	Velocity_Cache_3_4_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[95*3*DATA_WIDTH-1:94*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(6)
	)
	Velocity_Cache_3_4_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[96*3*DATA_WIDTH-1:95*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(5),
		.CELL_Z(1)
	)
	Velocity_Cache_3_5_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[97*3*DATA_WIDTH-1:96*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(5),
		.CELL_Z(2)
	)
	Velocity_Cache_3_5_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[98*3*DATA_WIDTH-1:97*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(5),
		.CELL_Z(3)
	)
	Velocity_Cache_3_5_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[99*3*DATA_WIDTH-1:98*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(5),
		.CELL_Z(4)
	)
	Velocity_Cache_3_5_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[100*3*DATA_WIDTH-1:99*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(5),
		.CELL_Z(5)
	)
	Velocity_Cache_3_5_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[101*3*DATA_WIDTH-1:100*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(5),
		.CELL_Z(6)
	)
	Velocity_Cache_3_5_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[102*3*DATA_WIDTH-1:101*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(6),
		.CELL_Z(1)
	)
	Velocity_Cache_3_6_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[103*3*DATA_WIDTH-1:102*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(6),
		.CELL_Z(2)
	)
	Velocity_Cache_3_6_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[104*3*DATA_WIDTH-1:103*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(6),
		.CELL_Z(3)
	)
	Velocity_Cache_3_6_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[105*3*DATA_WIDTH-1:104*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(6),
		.CELL_Z(4)
	)
	Velocity_Cache_3_6_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[106*3*DATA_WIDTH-1:105*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(6),
		.CELL_Z(5)
	)
	Velocity_Cache_3_6_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[107*3*DATA_WIDTH-1:106*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(6),
		.CELL_Z(6)
	)
	Velocity_Cache_3_6_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[108*3*DATA_WIDTH-1:107*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(1)
	)
	Velocity_Cache_4_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[109*3*DATA_WIDTH-1:108*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(2)
	)
	Velocity_Cache_4_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[110*3*DATA_WIDTH-1:109*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(3)
	)
	Velocity_Cache_4_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[111*3*DATA_WIDTH-1:110*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(4)
	)
	Velocity_Cache_4_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[112*3*DATA_WIDTH-1:111*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(5)
	)
	Velocity_Cache_4_1_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[113*3*DATA_WIDTH-1:112*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(6)
	)
	Velocity_Cache_4_1_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[114*3*DATA_WIDTH-1:113*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(1)
	)
	Velocity_Cache_4_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[115*3*DATA_WIDTH-1:114*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(2)
	)
	Velocity_Cache_4_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[116*3*DATA_WIDTH-1:115*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(3)
	)
	Velocity_Cache_4_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[117*3*DATA_WIDTH-1:116*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(4)
	)
	Velocity_Cache_4_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[118*3*DATA_WIDTH-1:117*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(5)
	)
	Velocity_Cache_4_2_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[119*3*DATA_WIDTH-1:118*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(6)
	)
	Velocity_Cache_4_2_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[120*3*DATA_WIDTH-1:119*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(1)
	)
	Velocity_Cache_4_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[121*3*DATA_WIDTH-1:120*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(2)
	)
	Velocity_Cache_4_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[122*3*DATA_WIDTH-1:121*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(3)
	)
	Velocity_Cache_4_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[123*3*DATA_WIDTH-1:122*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(4)
	)
	Velocity_Cache_4_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[124*3*DATA_WIDTH-1:123*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(5)
	)
	Velocity_Cache_4_3_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[125*3*DATA_WIDTH-1:124*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(6)
	)
	Velocity_Cache_4_3_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[126*3*DATA_WIDTH-1:125*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(1)
	)
	Velocity_Cache_4_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[127*3*DATA_WIDTH-1:126*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(2)
	)
	Velocity_Cache_4_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[128*3*DATA_WIDTH-1:127*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(3)
	)
	Velocity_Cache_4_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[129*3*DATA_WIDTH-1:128*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(4)
	)
	Velocity_Cache_4_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[130*3*DATA_WIDTH-1:129*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(5)
	)
	Velocity_Cache_4_4_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[131*3*DATA_WIDTH-1:130*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(6)
	)
	Velocity_Cache_4_4_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[132*3*DATA_WIDTH-1:131*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(5),
		.CELL_Z(1)
	)
	Velocity_Cache_4_5_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[133*3*DATA_WIDTH-1:132*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(5),
		.CELL_Z(2)
	)
	Velocity_Cache_4_5_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[134*3*DATA_WIDTH-1:133*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(5),
		.CELL_Z(3)
	)
	Velocity_Cache_4_5_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[135*3*DATA_WIDTH-1:134*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(5),
		.CELL_Z(4)
	)
	Velocity_Cache_4_5_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[136*3*DATA_WIDTH-1:135*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(5),
		.CELL_Z(5)
	)
	Velocity_Cache_4_5_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[137*3*DATA_WIDTH-1:136*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(5),
		.CELL_Z(6)
	)
	Velocity_Cache_4_5_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[138*3*DATA_WIDTH-1:137*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(6),
		.CELL_Z(1)
	)
	Velocity_Cache_4_6_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[139*3*DATA_WIDTH-1:138*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(6),
		.CELL_Z(2)
	)
	Velocity_Cache_4_6_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[140*3*DATA_WIDTH-1:139*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(6),
		.CELL_Z(3)
	)
	Velocity_Cache_4_6_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[141*3*DATA_WIDTH-1:140*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(6),
		.CELL_Z(4)
	)
	Velocity_Cache_4_6_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[142*3*DATA_WIDTH-1:141*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(6),
		.CELL_Z(5)
	)
	Velocity_Cache_4_6_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[143*3*DATA_WIDTH-1:142*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(6),
		.CELL_Z(6)
	)
	Velocity_Cache_4_6_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[144*3*DATA_WIDTH-1:143*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(1),
		.CELL_Z(1)
	)
	Velocity_Cache_5_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[145*3*DATA_WIDTH-1:144*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(1),
		.CELL_Z(2)
	)
	Velocity_Cache_5_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[146*3*DATA_WIDTH-1:145*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(1),
		.CELL_Z(3)
	)
	Velocity_Cache_5_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[147*3*DATA_WIDTH-1:146*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(1),
		.CELL_Z(4)
	)
	Velocity_Cache_5_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[148*3*DATA_WIDTH-1:147*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(1),
		.CELL_Z(5)
	)
	Velocity_Cache_5_1_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[149*3*DATA_WIDTH-1:148*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(1),
		.CELL_Z(6)
	)
	Velocity_Cache_5_1_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[150*3*DATA_WIDTH-1:149*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(2),
		.CELL_Z(1)
	)
	Velocity_Cache_5_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[151*3*DATA_WIDTH-1:150*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(2),
		.CELL_Z(2)
	)
	Velocity_Cache_5_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[152*3*DATA_WIDTH-1:151*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(2),
		.CELL_Z(3)
	)
	Velocity_Cache_5_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[153*3*DATA_WIDTH-1:152*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(2),
		.CELL_Z(4)
	)
	Velocity_Cache_5_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[154*3*DATA_WIDTH-1:153*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(2),
		.CELL_Z(5)
	)
	Velocity_Cache_5_2_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[155*3*DATA_WIDTH-1:154*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(2),
		.CELL_Z(6)
	)
	Velocity_Cache_5_2_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[156*3*DATA_WIDTH-1:155*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(3),
		.CELL_Z(1)
	)
	Velocity_Cache_5_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[157*3*DATA_WIDTH-1:156*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(3),
		.CELL_Z(2)
	)
	Velocity_Cache_5_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[158*3*DATA_WIDTH-1:157*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(3),
		.CELL_Z(3)
	)
	Velocity_Cache_5_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[159*3*DATA_WIDTH-1:158*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(3),
		.CELL_Z(4)
	)
	Velocity_Cache_5_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[160*3*DATA_WIDTH-1:159*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(3),
		.CELL_Z(5)
	)
	Velocity_Cache_5_3_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[161*3*DATA_WIDTH-1:160*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(3),
		.CELL_Z(6)
	)
	Velocity_Cache_5_3_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[162*3*DATA_WIDTH-1:161*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(4),
		.CELL_Z(1)
	)
	Velocity_Cache_5_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[163*3*DATA_WIDTH-1:162*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(4),
		.CELL_Z(2)
	)
	Velocity_Cache_5_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[164*3*DATA_WIDTH-1:163*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(4),
		.CELL_Z(3)
	)
	Velocity_Cache_5_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[165*3*DATA_WIDTH-1:164*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(4),
		.CELL_Z(4)
	)
	Velocity_Cache_5_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[166*3*DATA_WIDTH-1:165*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(4),
		.CELL_Z(5)
	)
	Velocity_Cache_5_4_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[167*3*DATA_WIDTH-1:166*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(4),
		.CELL_Z(6)
	)
	Velocity_Cache_5_4_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[168*3*DATA_WIDTH-1:167*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(5),
		.CELL_Z(1)
	)
	Velocity_Cache_5_5_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[169*3*DATA_WIDTH-1:168*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(5),
		.CELL_Z(2)
	)
	Velocity_Cache_5_5_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[170*3*DATA_WIDTH-1:169*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(5),
		.CELL_Z(3)
	)
	Velocity_Cache_5_5_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[171*3*DATA_WIDTH-1:170*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(5),
		.CELL_Z(4)
	)
	Velocity_Cache_5_5_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[172*3*DATA_WIDTH-1:171*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(5),
		.CELL_Z(5)
	)
	Velocity_Cache_5_5_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[173*3*DATA_WIDTH-1:172*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(5),
		.CELL_Z(6)
	)
	Velocity_Cache_5_5_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[174*3*DATA_WIDTH-1:173*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(6),
		.CELL_Z(1)
	)
	Velocity_Cache_5_6_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[175*3*DATA_WIDTH-1:174*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(6),
		.CELL_Z(2)
	)
	Velocity_Cache_5_6_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[176*3*DATA_WIDTH-1:175*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(6),
		.CELL_Z(3)
	)
	Velocity_Cache_5_6_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[177*3*DATA_WIDTH-1:176*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(6),
		.CELL_Z(4)
	)
	Velocity_Cache_5_6_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[178*3*DATA_WIDTH-1:177*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(6),
		.CELL_Z(5)
	)
	Velocity_Cache_5_6_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[179*3*DATA_WIDTH-1:178*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_Y(6),
		.CELL_Z(6)
	)
	Velocity_Cache_5_6_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[180*3*DATA_WIDTH-1:179*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(1),
		.CELL_Z(1)
	)
	Velocity_Cache_6_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[181*3*DATA_WIDTH-1:180*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(1),
		.CELL_Z(2)
	)
	Velocity_Cache_6_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[182*3*DATA_WIDTH-1:181*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(1),
		.CELL_Z(3)
	)
	Velocity_Cache_6_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[183*3*DATA_WIDTH-1:182*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(1),
		.CELL_Z(4)
	)
	Velocity_Cache_6_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[184*3*DATA_WIDTH-1:183*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(1),
		.CELL_Z(5)
	)
	Velocity_Cache_6_1_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[185*3*DATA_WIDTH-1:184*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(1),
		.CELL_Z(6)
	)
	Velocity_Cache_6_1_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[186*3*DATA_WIDTH-1:185*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(2),
		.CELL_Z(1)
	)
	Velocity_Cache_6_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[187*3*DATA_WIDTH-1:186*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(2),
		.CELL_Z(2)
	)
	Velocity_Cache_6_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[188*3*DATA_WIDTH-1:187*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(2),
		.CELL_Z(3)
	)
	Velocity_Cache_6_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[189*3*DATA_WIDTH-1:188*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(2),
		.CELL_Z(4)
	)
	Velocity_Cache_6_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[190*3*DATA_WIDTH-1:189*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(2),
		.CELL_Z(5)
	)
	Velocity_Cache_6_2_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[191*3*DATA_WIDTH-1:190*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(2),
		.CELL_Z(6)
	)
	Velocity_Cache_6_2_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[192*3*DATA_WIDTH-1:191*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(3),
		.CELL_Z(1)
	)
	Velocity_Cache_6_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[193*3*DATA_WIDTH-1:192*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(3),
		.CELL_Z(2)
	)
	Velocity_Cache_6_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[194*3*DATA_WIDTH-1:193*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(3),
		.CELL_Z(3)
	)
	Velocity_Cache_6_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[195*3*DATA_WIDTH-1:194*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(3),
		.CELL_Z(4)
	)
	Velocity_Cache_6_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[196*3*DATA_WIDTH-1:195*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(3),
		.CELL_Z(5)
	)
	Velocity_Cache_6_3_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[197*3*DATA_WIDTH-1:196*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(3),
		.CELL_Z(6)
	)
	Velocity_Cache_6_3_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[198*3*DATA_WIDTH-1:197*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(4),
		.CELL_Z(1)
	)
	Velocity_Cache_6_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[199*3*DATA_WIDTH-1:198*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(4),
		.CELL_Z(2)
	)
	Velocity_Cache_6_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[200*3*DATA_WIDTH-1:199*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(4),
		.CELL_Z(3)
	)
	Velocity_Cache_6_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[201*3*DATA_WIDTH-1:200*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(4),
		.CELL_Z(4)
	)
	Velocity_Cache_6_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[202*3*DATA_WIDTH-1:201*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(4),
		.CELL_Z(5)
	)
	Velocity_Cache_6_4_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[203*3*DATA_WIDTH-1:202*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(4),
		.CELL_Z(6)
	)
	Velocity_Cache_6_4_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[204*3*DATA_WIDTH-1:203*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(5),
		.CELL_Z(1)
	)
	Velocity_Cache_6_5_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[205*3*DATA_WIDTH-1:204*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(5),
		.CELL_Z(2)
	)
	Velocity_Cache_6_5_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[206*3*DATA_WIDTH-1:205*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(5),
		.CELL_Z(3)
	)
	Velocity_Cache_6_5_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[207*3*DATA_WIDTH-1:206*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(5),
		.CELL_Z(4)
	)
	Velocity_Cache_6_5_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[208*3*DATA_WIDTH-1:207*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(5),
		.CELL_Z(5)
	)
	Velocity_Cache_6_5_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[209*3*DATA_WIDTH-1:208*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(5),
		.CELL_Z(6)
	)
	Velocity_Cache_6_5_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[210*3*DATA_WIDTH-1:209*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(6),
		.CELL_Z(1)
	)
	Velocity_Cache_6_6_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[211*3*DATA_WIDTH-1:210*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(6),
		.CELL_Z(2)
	)
	Velocity_Cache_6_6_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[212*3*DATA_WIDTH-1:211*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(6),
		.CELL_Z(3)
	)
	Velocity_Cache_6_6_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[213*3*DATA_WIDTH-1:212*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(6),
		.CELL_Z(4)
	)
	Velocity_Cache_6_6_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[214*3*DATA_WIDTH-1:213*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(6),
		.CELL_Z(5)
	)
	Velocity_Cache_6_6_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[215*3*DATA_WIDTH-1:214*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(6),
		.CELL_Y(6),
		.CELL_Z(6)
	)
	Velocity_Cache_6_6_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[216*3*DATA_WIDTH-1:215*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(1),
		.CELL_Z(1)
	)
	Velocity_Cache_7_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[217*3*DATA_WIDTH-1:216*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(1),
		.CELL_Z(2)
	)
	Velocity_Cache_7_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[218*3*DATA_WIDTH-1:217*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(1),
		.CELL_Z(3)
	)
	Velocity_Cache_7_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[219*3*DATA_WIDTH-1:218*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(1),
		.CELL_Z(4)
	)
	Velocity_Cache_7_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[220*3*DATA_WIDTH-1:219*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(1),
		.CELL_Z(5)
	)
	Velocity_Cache_7_1_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[221*3*DATA_WIDTH-1:220*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(1),
		.CELL_Z(6)
	)
	Velocity_Cache_7_1_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[222*3*DATA_WIDTH-1:221*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(2),
		.CELL_Z(1)
	)
	Velocity_Cache_7_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[223*3*DATA_WIDTH-1:222*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(2),
		.CELL_Z(2)
	)
	Velocity_Cache_7_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[224*3*DATA_WIDTH-1:223*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(2),
		.CELL_Z(3)
	)
	Velocity_Cache_7_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[225*3*DATA_WIDTH-1:224*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(2),
		.CELL_Z(4)
	)
	Velocity_Cache_7_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[226*3*DATA_WIDTH-1:225*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(2),
		.CELL_Z(5)
	)
	Velocity_Cache_7_2_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[227*3*DATA_WIDTH-1:226*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(2),
		.CELL_Z(6)
	)
	Velocity_Cache_7_2_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[228*3*DATA_WIDTH-1:227*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(3),
		.CELL_Z(1)
	)
	Velocity_Cache_7_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[229*3*DATA_WIDTH-1:228*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(3),
		.CELL_Z(2)
	)
	Velocity_Cache_7_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[230*3*DATA_WIDTH-1:229*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(3),
		.CELL_Z(3)
	)
	Velocity_Cache_7_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[231*3*DATA_WIDTH-1:230*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(3),
		.CELL_Z(4)
	)
	Velocity_Cache_7_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[232*3*DATA_WIDTH-1:231*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(3),
		.CELL_Z(5)
	)
	Velocity_Cache_7_3_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[233*3*DATA_WIDTH-1:232*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(3),
		.CELL_Z(6)
	)
	Velocity_Cache_7_3_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[234*3*DATA_WIDTH-1:233*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(4),
		.CELL_Z(1)
	)
	Velocity_Cache_7_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[235*3*DATA_WIDTH-1:234*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(4),
		.CELL_Z(2)
	)
	Velocity_Cache_7_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[236*3*DATA_WIDTH-1:235*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(4),
		.CELL_Z(3)
	)
	Velocity_Cache_7_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[237*3*DATA_WIDTH-1:236*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(4),
		.CELL_Z(4)
	)
	Velocity_Cache_7_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[238*3*DATA_WIDTH-1:237*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(4),
		.CELL_Z(5)
	)
	Velocity_Cache_7_4_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[239*3*DATA_WIDTH-1:238*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(4),
		.CELL_Z(6)
	)
	Velocity_Cache_7_4_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[240*3*DATA_WIDTH-1:239*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(5),
		.CELL_Z(1)
	)
	Velocity_Cache_7_5_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[241*3*DATA_WIDTH-1:240*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(5),
		.CELL_Z(2)
	)
	Velocity_Cache_7_5_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[242*3*DATA_WIDTH-1:241*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(5),
		.CELL_Z(3)
	)
	Velocity_Cache_7_5_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[243*3*DATA_WIDTH-1:242*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(5),
		.CELL_Z(4)
	)
	Velocity_Cache_7_5_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[244*3*DATA_WIDTH-1:243*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(5),
		.CELL_Z(5)
	)
	Velocity_Cache_7_5_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[245*3*DATA_WIDTH-1:244*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(5),
		.CELL_Z(6)
	)
	Velocity_Cache_7_5_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[246*3*DATA_WIDTH-1:245*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(6),
		.CELL_Z(1)
	)
	Velocity_Cache_7_6_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[247*3*DATA_WIDTH-1:246*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(6),
		.CELL_Z(2)
	)
	Velocity_Cache_7_6_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[248*3*DATA_WIDTH-1:247*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(6),
		.CELL_Z(3)
	)
	Velocity_Cache_7_6_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[249*3*DATA_WIDTH-1:248*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(6),
		.CELL_Z(4)
	)
	Velocity_Cache_7_6_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[250*3*DATA_WIDTH-1:249*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(6),
		.CELL_Z(5)
	)
	Velocity_Cache_7_6_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[251*3*DATA_WIDTH-1:250*3*DATA_WIDTH])
	);

	Velocity_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),									// Data width of a single force value, 32-bit
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(7),
		.CELL_Y(6),
		.CELL_Z(6)
	)
	Velocity_Cache_7_6_6
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_velocity_read_addr),
		.in_data(Motion_Update_out_velocity_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_velocity_data_valid),		// Signify if the new incoming data is valid
		.in_rden(Motion_Update_velocity_read_en),
		.out_particle_info(wire_cache_to_motion_update_velocity_data[252*3*DATA_WIDTH-1:251*3*DATA_WIDTH])
	);

endmodule
